���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.5.2�ub�n_estimators�K�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��numpy._core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��ExerciseAngina��Oldpeak��ST_Slope�et�b�n_features_in_�K�
_n_samples�M��
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�_n_samples_bootstrap�M��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ�
hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��h3�f8�����R�(KhQNNNJ����J����K t�b�C              �?�t�bhUh'�scalar���hPC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hK�
node_count�K��nodes�h)h,K ��h.��R�(KK���h3�V64�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h�hPK ��h�hPK��h�hPK��h�hbK��h�hbK ��h�hPK(��h�hbK0��h�h3�u1�����R�(Kh7NNNJ����J����K t�bK8��uK@KKt�b�B@0         b                    @j8je3�?�           ��@                                   �?"\�����?�             t@                      
             �?���W���?8            �U@                                   �?$��m��?             :@                                 �u@�GN�z�?             6@                                  �?�����H�?             2@                                  �?z�G�z�?             $@              	                   �n@�����H�?             "@        ������������������������       �                     @        
                          �p@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                  �}@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        (             N@               1       	             �?��Q:��?�            �m@                                 �X@�ӭ�a��?a             b@                                   @I@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @               &                   pq@��)��g�?[             a@                                  �?4�0_���?J            @\@                                  �`@���Q��?             @        ������������������������       �                     �?                                  �d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                %       
             �?��Wv��?F             [@        !       "       
             �?��
ц��?             *@        ������������������������       �                     @        #       $                   0f@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        ;            �W@        '       (                    @E@�q�q�?             8@        ������������������������       �                     (@        )       *                   �`@�q�q�?
             (@        ������������������������       �                     �?        +       ,       
             �?���|���?	             &@        ������������������������       �                     @        -       .                   �q@�q�q�?             @        ������������������������       �                     �?        /       0                    �N@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        2       W       
             �?���j��?7             W@       3       8                    �F@6��f�?+            @S@        4       7                    �?�q�q�?             @        5       6       	              @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        9       H                   �h@�ˡ�5��?%            �Q@        :       A       	          033�?��X��?             <@       ;       @       	          ����?��.k���?	             1@       <       =                   @`@�	j*D�?             *@       ������������������������       �                     @        >       ?                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        B       C                    �?�C��2(�?             &@        ������������������������       �                     @        D       E       
             �?z�G�z�?             @        ������������������������       �                     @        F       G                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       J                    @N@Du9iH��?            �E@        ������������������������       �                     :@        K       P                    �?@�0�!��?             1@        L       O       	          ���@���Q��?             @       M       N                    �P@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        Q       V                    �?�8��8��?             (@       R       U                   m@r�q��?             @        S       T                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        X       Y                   `U@�q�q�?             .@        ������������������������       �                      @        Z       [                   Pi@�θ�?
             *@        ������������������������       �                     @        \       _                    �?      �?              @       ]       ^                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        `       a                   �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        c       �                    �?�}�	���?           �y@       d       �                   �e@�������?�            �s@       e       �       
             �?H.�!���?�            �r@       f       �                   pn@L�'�7��?�            @m@       g       l                   �g@`	�<��?T            �a@        h       i                   @a@ _�@�Y�?#             M@       ������������������������       �                     J@        j       k                    @J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        m       t                   0j@�?a/��?1            �T@        n       s                   �i@���|���?             6@       o       r       	          ����?�d�����?             3@        p       q       	          ����?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        u       �       	          ����?��.��?#            �N@        v       y       	             �?      �?             4@        w       x                    m@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        z                           �?�����H�?             "@       {       |                    �?r�q��?             @        ������������������������       �                      @        }       ~                   pm@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        �       �                   q@�g�y��?:            @W@        ������������������������       �                    �B@        �       �                    �?�h����?#             L@        ������������������������       �        
             4@        �       �                    �?�8��8��?             B@       �       �                     M@r�q��?             2@       �       �       	          ����?$�q-�?
             *@        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �       	             �?���Q��?             @        ������������������������       �                     �?        �       �                   0r@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     2@        �       �                    �?�q�q�?0            �P@       �       �                   �_@��x_F-�?$            �I@       �       �       	          ����?�n_Y�K�?             :@       �       �       	          ����?z�G�z�?             4@       �       �                   0e@@�0�!��?             1@       �       �                   �b@��S�ۿ?             .@       ������������������������       �                     $@        �       �                   �c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    ]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     9@        �       �                    c@z�G�z�?             .@       �       �       	          ����?؇���X�?             ,@       ������������������������       �                      @        �       �                   ``@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?$�q-�?             *@        �       �                   l@      �?             @       �       �                    h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �       
             �?�FVQ&�?=            �X@       �       �                   Pz@XB���?4            �U@       �       �                    �R@ ��N8�?2             U@       ������������������������       �        0            �T@        �       �                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   ��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    Z@      �?	             (@        ������������������������       �                     �?        �       �                    �?"pc�
�?             &@       ������������������������       �                     @        �       �                    @K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �t�b�values�h)h,K ��h.��R�(KK�KK��hb�B  ���Y��?t�S��?.>9\�?ǣ���G�?*kʚ���?���)kʺ?�N��N��?vb'vb'�?�袋.��?]t�E�?�q�q�?�q�q�?�������?�������?�q�q�?�q�q�?      �?        �������?�������?              �?      �?                      �?      �?              �?      �?              �?      �?                      �?      �?        'u_[�?�A�I��?�q�q�?�8��8��?�$I�$I�?۶m۶m�?      �?                      �?/�#EC�?������?�8�1�s�?�:Fq�c�?333333�?�������?              �?      �?      �?      �?                      �?�^B{	��?{	�%���?�؉�؉�?�;�;�?      �?              �?      �?              �?      �?              �?        �������?�������?      �?        �������?�������?      �?        F]t�E�?]t�E]�?              �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?!Y�B�?ozӛ���?�cj`��?g�'�Y�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        H���@��?�RO�o��?%I�$I��?n۶m۶�?�?�������?;�;��?vb'vb'�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        F]t�E�?]t�E�?              �?�������?�������?              �?      �?      �?              �?      �?        w�qGܱ?qG�w��?              �?�������?ZZZZZZ�?�������?333333�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?ى�؉��?�؉�؉�?      �?              �?      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ����?��R�y�?�:x����?G�
��?)\���(�?�(\����?���?�������?E�)͋?�?o����?�{a���?#,�4�r�?              �?UUUUUU�?�������?              �?      �?        rY1P��?x���k�?F]t�E�?]t�E]�?y�5���?Cy�5��?r�q��?�q�q�?              �?      �?                      �?      �?        ������?�����?      �?      �?F]t�E�?/�袋.�?              �?      �?        �q�q�?�q�q�?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?�B!��?��{���?              �?۶m۶m�?�$I�$I�?              �?UUUUUU�?UUUUUU�?UUUUUU�?�������?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?333333�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?�������?�?;�;��?ى�؉��?�������?�������?ZZZZZZ�?�������?�������?�?      �?        �������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?�������?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �؉�؉�?;�;��?      �?      �?      �?      �?      �?                      �?      �?              �?        |���?>����?�{a���?GX�i���?�a�a�?�y��y��?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?        F]t�E�?/�袋.�?              �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ/��hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@/         l       
             �?4�5����?�           ��@              /                    @P� �&�?           @y@                                   �?���e��?X            �`@                                  �g@�>4և��?             <@                                   �G@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @               	                    �I@���}<S�?             7@        ������������������������       �                     $@        
                           �?8�Z$���?             *@       ������������������������       �        	             &@        ������������������������       �                      @                                  0i@�3�E���?D             Z@                                  �c@������?            �B@       ������������������������       �                     ?@                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                   �b@�#}7��?.            �P@                                 �\@z�G�z�?             D@                                  @m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                      	          ����?$G$n��?            �B@                                  �]@     ��?             0@        ������������������������       �                     @                                  @e@      �?             $@                                 Pa@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     5@        !       "                   �l@�5��?             ;@        ������������������������       �                      @        #       *                    �?D�n�3�?             3@       $       '                    �?�q�q�?             "@       %       &       	             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        (       )                   pf@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        +       .                   �b@      �?             $@       ,       -                   `m@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        0       1       	          ����?l��\��?�             q@        ������������������������       �                    �I@        2       9                   `[@H �/$��?�            �k@        3       4       	          hff�?      �?"             P@        ������������������������       �                     �?        5       8                   �Q@ ������?!            �O@        6       7                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �N@        :       G                    �?��V���?j            �c@        ;       F       	          ����?���|���?            �@@       <       E                    �O@�eP*L��?             6@       =       >                    @D@      �?	             0@        ������������������������       �                      @        ?       @                   @m@؇���X�?             ,@        ������������������������       �                     @        A       D                    �M@      �?              @       B       C                   @`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        H       I                   �U@6uH���?W             _@        ������������������������       �                     �?        J       U                    \@��p\�?V            �^@        K       L                   @Z@������?
             1@        ������������������������       �                     @        M       T                    �M@���Q��?             $@       N       S                   p@և���X�?             @       O       R                    �I@z�G�z�?             @       P       Q                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        V       ]       	          ����?����?L            �Z@        W       Z       	          ����?����X�?             @        X       Y                    X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        [       \                   �`@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ^       k                    �R@Pa�	�?G            �X@       _       f                    �?@�E�x�?F            �X@        `       a       	          033�?�8��8��?
             (@        ������������������������       �                     @        b       e       	             �?r�q��?             @        c       d                    @P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        g       j                   �_@��f�{��?<            �U@        h       i                    \@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �        
             ,@        ������������������������       �        1            �Q@        ������������������������       �                     �?        m       |                   @E@`}�?��?�            �t@        n       {                    �?P����?             C@        o       v                    �K@��Q��?             4@        p       q                    ]@      �?              @        ������������������������       �                      @        r       s                    @r�q��?             @        ������������������������       �                      @        t       u                   @_@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        w       x                    `P@r�q��?             (@       ������������������������       �                     @        y       z                    `R@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        }       �                    @L@�@i����?�            @r@       ~                           �?�uR����?�            �k@        ������������������������       �        $            �P@        �       �       	          033�?�Z��=��?b            �c@       �       �                    @�H��Ԉ�?]            �b@       �       �                    �?�&=�w��?B            �Z@       �       �                   @[@�E�����?:            �V@        �       �                   @Y@�q�q�?             @        ������������������������       �                     �?        �       �                    @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        7            �U@        �       �                   �g@     ��?             0@       ������������������������       �                     (@        �       �                   �h@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �b@�<ݚ�?            �F@       ������������������������       �                     9@        �       �                   �f@      �?             4@       �       �                    �?�q�q�?
             .@       �       �       	             �?      �?             $@       �       �                   �e@�q�q�?             @       �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��x�5��?*            @Q@       �       �                    �M@�\�u��?            �I@        �       �                    d@      �?             6@       �       �                   �b@����X�?	             ,@       �       �                   Hp@"pc�
�?             &@       ������������������������       �                      @        �       �                   0b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    \@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          033@д>��C�?             =@       �       �                    �O@؇���X�?             <@        ������������������������       �                     .@        �       �                     P@�	j*D�?
             *@        ������������������������       �                      @        �       �                    @"pc�
�?	             &@       ������������������������       �                     @        �       �                    ]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�q�q�?             2@        ������������������������       �                     @        ������������������������       �                     (@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�   Np	�?���Gw{�?
L:5r�?�l�2|#�?>���>�?�>���?�$I�$I�?�m۶m��?�������?333333�?      �?                      �?ӛ���7�?d!Y�B�?      �?        ;�;��?;�;��?      �?                      �?ى�؉��?;�;��?к����?��g�`��?              �?UUUUUU�?UUUUUU�?              �?      �?        ���[��?~5&��?ffffff�?ffffff�?UUUUUU�?UUUUUU�?      �?                      �?���L�?к����?      �?      �?              �?      �?      �?      �?      �?      �?                      �?              �?              �?h/�����?/�����?      �?        (������?l(�����?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?              �?      �?                      �?�������?------�?              �?�ͻ?�^��^��?      �?      �?      �?        AA�?��}��}�?      �?      �?              �?      �?                      �?������?����?F]t�E�?]t�E]�?t�E]t�?]t�E�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?      �?                      �?      �?                      �?              �?��RJ)��?k���Zk�?      �?        ��+Q��?�]�ڕ��?�?xxxxxx�?              �?�������?333333�?�$I�$I�?۶m۶m�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?�V�9�&�?��`��}�?�$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?              �?      �?        |���?|���?9/���?և���X�?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�}A_Ї?������?�?�������?      �?                      �?              �?      �?        �בz�?�[����?Q^Cy��?�P^Cy�?�������?ffffff�?      �?      �?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?        �������?UUUUUU�?      �?        333333�?�������?              �?      �?                      �?X�^�z��?�B�
*�?V�-(�j�?O���橴?      �?        t��0�T�?b��x�Y�?�!�z�?��^x/��?tHM0���?�x+�R�?P��O���?l�l��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?      �?      �?              �?      �?              �?      �?        9��8���?�q�q�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?      �?      �?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?0�̵�?�Q�g���?�������?�?      �?      �?�m۶m��?�$I�$I�?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?a���{�?|a���?۶m۶m�?�$I�$I�?      �?        vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?      �?              �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJu�7hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKɅ�h��B@2         J       	          ����?p�Vv���?�           ��@               3                    �?X~�pX��?�            �v@                     
             �?BA�V�?�            �r@               	                    �?      �?0             R@                                  �Q@      �?	             (@        ������������������������       �                      @                                   @ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        
              	          833�?R���Q�?'             N@                                 `c@p���?             I@       ������������������������       �                    �F@                                  �d@z�G�z�?             @                                  �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?z�G�z�?             $@                                 q@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                    @ d�=��?�            @l@                                 Hp@PA��ڡ?k             e@       ������������������������       �        R            �`@                                  Xp@l��\��?             A@        ������������������������       �                      @                                  pq@      �?             @@        ������������������������       �        
             0@                                  �g@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        !       "       	             ࿜MWl��?#            �L@        ������������������������       �                     �?        #       $                    P@d}h���?"             L@        ������������������������       �                     @        %       0                    �M@8�Z$���?             J@       &       /                   l@��(\���?             D@       '       ,                    �?�LQ�1	�?             7@       (       +                    �D@�KM�]�?
             3@        )       *                    a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        -       .                     G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        1       2                   �b@�q�q�?             (@       ������������������������       �                     @        ������������������������       �                     @        4       I                   Pd@��y�:�?,            �P@       5       8                    [@^l��[B�?'             M@        6       7                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        9       >                   �n@�+$�jP�?$             K@       :       ;                   �`@      �?             @@       ������������������������       �                     :@        <       =                    b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       D                     N@8�A�0��?             6@        @       A                    �?"pc�
�?             &@       ������������������������       �                     @        B       C                   �b@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        E       F                   `Y@���|���?             &@        ������������������������       �                      @        G       H                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        K       �       	          033�?�zц��?�            w@        L       c                    @���m�?]             b@        M       R                    �?�"U����?             �I@        N       Q                    �?      �?
             0@        O       P       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        S       b                    �N@��
P��?            �A@       T       U                   �[@`�Q��?             9@        ������������������������       �                     @        V       Y                    _@��s����?             5@        W       X                    @M@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        Z       [                   �`@�����H�?
             2@        ������������������������       �                      @        \       ]                    @K@z�G�z�?             $@        ������������������������       �                     @        ^       _                    �?      �?             @        ������������������������       �                     �?        `       a                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        d       k                   �X@��E�B��?=            �W@        e       j                   �`@��
ц��?             *@       f       g                   �Y@      �?              @        ������������������������       �                     �?        h       i                   @\@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        l       {                   pb@�>����?6            @T@       m       p                   �[@hA� �?.            �Q@        n       o                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        q       r                   pa@Pa�	�?,            �P@       ������������������������       �                    �C@        s       z                   �u@�>����?             ;@       t       y                   �a@ ��WV�?             :@        u       v                    �?z�G�z�?             @        ������������������������       �                      @        w       x       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        ������������������������       �                     �?        |       �                     L@���!pc�?             &@        }       �                    �J@      �?             @       ~       �                    �?      �?             @              �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?������?�             l@        �       �       
             �?��
P�?3            �Q@       �       �                   `_@ {��e�?&            �J@        �       �                    @O@�q�q�?             2@       ������������������������       �                     &@        �       �       	             @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   d@؇���X�?            �A@       �       �                    �?ףp=
�?             >@       �       �       	          `ff�?z�G�z�?             .@        �       �                   �\@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �       	          ���@r�q��?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        �       �                   pe@���Q��?             @       �       �                    �L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     Q@��.k���?             1@       �       �                   @b@���Q��?             .@       �       �                    �?"pc�
�?	             &@       �       �                    �?�q�q�?             @       �       �                     I@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   8q@@4և���?e            @c@       �       �                    Z@t��%�?N            �\@        �       �       	             @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @��X��?L             \@        �       �                   �a@d}h���?             ,@       �       �                    �J@      �?              @        �       �                   �l@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   0c@��<D�m�?A            �X@       �       �       	          ����?hl �&�?>             W@        �       �                    @L@�C��2(�?             6@       ������������������������       �        	             .@        �       �                   @^@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       	          033@`����֜?/            �Q@       ������������������������       �        !            �H@        �       �                   �_@���N8�?             5@        �       �       	          `ff
@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        �       �                   �p@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �C@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  w
��,@�?�z�����?�^�z���?�B�
*�?�Ug�{�?`��c.�?      �?      �?      �?      �?              �?�������?�������?      �?                      �?333333�?333333�?{�G�z�?\���(\�?              �?�������?�������?      �?      �?              �?      �?                      �?�������?�������?�q�q�?�q�q�?      �?                      �?              �?���	��?x�!���?��s�n�?&�q-�?      �?        ------�?�������?              �?      �?      �?      �?              �?      �?      �?                      �?:��,���?�YLg1�?              �?I�$I�$�?۶m۶m�?              �?;�;��?;�;��?�������?333333�?��Moz��?Y�B��?�k(���?(�����?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?              �?        �������?�������?      �?                      �?~5&��?�@��~�?��=���?�=�����?      �?      �?      �?                      �?B{	�%��?/�����?      �?      �?              �?UUUUUU�?�������?              �?      �?        /�袋.�?颋.���?F]t�E�?/�袋.�?              �?�������?333333�?              �?      �?        ]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?                      �?      �?        o`E\��?@��(��?%�6Q�k�?m�d�&J�?�?�������?      �?      �?      �?      �?              �?      �?              �?        _�_��?PuPu�?��(\���?{�G�z�?              �?z��y���?�a�a�?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?      �?        �������?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?AL� &W�?�l�w6��?�؉�؉�?�;�;�?      �?      �?              �?۶m۶m�?�$I�$I�?              �?      �?                      �?h/�����?�Kh/��?_�_�?���?      �?      �?      �?                      �?|���?|���?              �?h/�����?�Kh/��?;�;��?O��N���?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        t�E]t�?F]t�E�?      �?      �?      �?      �?      �?      �?      �?                      �?              �?      �?                      �?I�$I�$�?n۶m۶�?�_�_�?uPuP�?
�[���?~�	�[�?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?                      �?�$I�$I�?۶m۶m�?�������?�������?�������?�������?�������?333333�?              �?      �?        �������?�������?              �?UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�?�������?�������?333333�?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?              �?              �?      �?              �?        �$I�$I�?n۶m۶�?�q�.�|�?�(�j��?UUUUUU�?UUUUUU�?              �?      �?        %I�$I��?۶m۶m�?۶m۶m�?I�$I�$�?      �?      �?      �?      �?      �?                      �?              �?              �?և���X�?��S�r
�?Y�B��?ozӛ���?F]t�E�?]t�E�?              �?�$I�$I�?�m۶m��?              �?      �?        �A�A�?�������?              �?�a�a�?��y��y�?      �?      �?      �?                      �?              �?      �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��!XhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKׅ�h��B�5         p                    �?U�ք�?�           ��@              [                    �?n�����?           @z@              ,       
             �?do@I�l�?�            �t@                                  �l@^H���+�?L            �[@              
       	          ����?X�<ݚ�?(             K@               	                     F@P���Q�?             4@                                    D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@                                   �?�!���?             A@        ������������������������       �                      @                      	          ����?
j*D>�?             :@        ������������������������       �                     "@                                  �c@ҳ�wY;�?             1@                                  @O@������?             .@       ������������������������       �                     "@                                  �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @               +                   �b@�d�����?$            �L@                                  �?~���L0�?!            �H@                                   �?�C��2(�?             &@                                  @_@      �?             @        ������������������������       �                      @                                  `X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               "       
             �?�?�'�@�?             C@                !                   e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        #       *                   0f@�#-���?            �A@       $       %                   �`@Pa�	�?            �@@       ������������������������       �                     8@        &       )                   0a@�����H�?             "@        '       (                   �n@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        -       J                    �?      �?�             l@       .       /                    �?�F�l���?            �g@        ������������������������       �        <            �V@        0       G                   ht@D���ͫ�?C            @Y@       1       B       	          ����?      �??             X@       2       5                   @E@X;��?;            @V@        3       4                    ^@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        6       A                   l@�Ń��̧?7             U@       7       >                    f@`�q�0ܴ?            �G@       8       9                    �?`���i��?             F@        ������������������������       �                      @        :       ;                    b@������?             B@       ������������������������       �                    �@@        <       =                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ?       @                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �B@        C       F                   �j@և���X�?             @       D       E                   0f@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        H       I                    �N@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        K       Z       	          833@"pc�
�?            �@@       L       U                    @     ��?             @@       M       N                    �?�>����?             ;@        ������������������������       �                     �?        O       P                    �? ��WV�?             :@        ������������������������       �                     @        Q       R                    �H@�}�+r��?             3@        ������������������������       �                     $@        S       T                   �e@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        V       Y                    p@���Q��?             @        W       X                   �f@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        \       g                    @M@ܻ�yX7�?4            @U@       ]       b                    @�q�q�?             H@        ^       a       
             �?���y4F�?             3@        _       `                   �a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        c       f       
             �?XB���?             =@        d       e                   �l@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     9@        h       m       
             �?�L���?            �B@       i       j                   `c@      �?             @@       ������������������������       �                     >@        k       l                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        n       o       	          ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        q       �       
             �?JN�#:�?�            �s@       r       �                    @pH����?�            �p@        s       |                   �`@�<ݚ�?&             K@       t       u                    �?��?^�k�?            �A@        ������������������������       �                      @        v       {                     N@ 7���B�?             ;@       w       x                    @M@��S�ۿ?
             .@       ������������������������       �                     &@        y       z       	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             (@        }       �       	             @D�n�3�?             3@       ~                          @_@ҳ�wY;�?             1@        ������������������������       �                     @        �       �       	          ����?      �?	             (@        ������������������������       �                     @        �       �       	          ����?�q�q�?             "@       �       �                   �a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   0a@��8����?�            �j@       �       �                    \@ ,U,?��?h            �d@        �       �                   �`@�Z��L��?,            �Q@        �       �                   @[@���y4F�?             3@       �       �       
             �?      �?             0@        ������������������������       �                      @        �       �                   `^@      �?              @        ������������������������       �                     @        �       �                   �Y@      �?             @        ������������������������       �                     �?        �       �                    Y@�q�q�?             @       �       �                   0j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?$�q-�?             J@       �       �       	             �?<���D�?            �@@       �       �                   `[@�X�<ݺ?             2@       ������������������������       �        
             1@        ������������������������       �                     �?        �       �                    �Q@z�G�z�?	             .@       ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     3@        �       �                    @L@ r���?<            �W@       ������������������������       �        !             J@        �       �                    �? �#�Ѵ�?            �E@       �       �                    �?      �?             @@        �       �                   `^@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `]@ 7���B�?             ;@        �       �                    Y@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     8@        ������������������������       �                     &@        �       �                   �m@      �?             H@       �       �       	             �?�+e�X�?             9@        �       �                    b@X�Cc�?             ,@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   �j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    \@�C��2(�?	             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     7@        �       �                    I@\X��t�?             G@        �       �                   b@�C��2(�?             &@       ������������������������       �                     "@        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?����X�?            �A@        ������������������������       �                     @        �       �                   ``@�q�q�?             >@        �       �                   @`@      �?	             ,@        ������������������������       �                     @        �       �                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @     ��?             0@        ������������������������       �                     @        �       �                    �?�z�G��?             $@       �       �                    �?և���X�?             @       �       �                   �b@���Q��?             @        ������������������������       �                     �?        �       �                    a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  ᓔ��?�5�;��?�Fk�Fk�?�r)�r)�?�N�����?�bѲ
n�?�g�`�|�?L�Ϻ��?�q�q�?r�q��?�������?ffffff�?�������?�������?              �?      �?                      �?�������?�������?      �?        b'vb'v�?;�;��?      �?        �������?�������?�?wwwwww�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        y�5���?Cy�5��?������?����>4�?]t�E�?F]t�E�?      �?      �?      �?              �?      �?              �?      �?              �?        y�5���?������?UUUUUU�?UUUUUU�?              �?      �?        _�_�?�A�A�?|���?|���?              �?�q�q�?�q�q�?      �?      �?      �?                      �?              �?      �?                      �?      �?      �?L�:,��?:kP<�q�?      �?        ��S� w�?��be�F�?      �?      �?�u�{���?�E(B�?�������?�������?      �?                      �?��<��<�?�a�a�?��F}g��?W�+�ɥ?F]t�E�?F]t�E�?      �?        �q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?333333�?�������?      �?                      �?/�袋.�?F]t�E�?      �?      �?�Kh/��?h/�����?              �?O��N���?;�;��?      �?        �5��P�?(�����?      �?        �q�q�?�q�q�?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�������?UUUUUU�?UUUUUU�?6��P^C�?(������?�������?�������?              �?      �?              �?        �{a���?GX�i���?      �?      �?              �?      �?                      �?L�Ϻ��?}���g�?      �?      �?              �?      �?      �?      �?                      �?�������?333333�?      �?                      �?I/�B�?.4`I/�?z�rv��?�1���?�q�q�?9��8���?�A�A�?_�_��?              �?h/�����?	�%����?�?�������?              �?      �?      �?      �?                      �?              �?l(�����?(������?�������?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?      �?      �?                      �?              �?�+J�#�?蝺����?��FS�׮?��ˊ��?��Vؼ?���.�d�?(������?6��P^C�?      �?      �?              �?      �?      �?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ;�;��?�؉�؉�?|���?|���?�q�q�?��8��8�?              �?      �?        �������?�������?              �?      �?                      �?�X�0Ҏ�?9�{n�S�?              �?�}A_Ч?�/����?      �?      �?�������?�������?      �?                      �?h/�����?	�%����?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?���Q��?R���Q�?�m۶m��?%I�$I��?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?]t�E�?      �?                      �?              �?!Y�B�?��Moz��?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?                      �?      �?      �?      �?        ffffff�?333333�?�$I�$I�?۶m۶m�?�������?333333�?      �?              �?      �?      �?                      �?      �?              �?        �t�bub�g     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJC�NhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@?         j                    @4�5����?�           ��@               U                    �?������?�            �t@              2                    @L@X�@��l�?�            �p@                     
             �?< 
2��?�            `i@                                  0a@\X��t�?             G@                                 pb@�q�q�?            �C@                      	              @�z�G��?             $@                     	          `ff�?և���X�?             @       	                           a@z�G�z�?             @       
                           �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                  �p@V�a�� �?             =@                     	             @����X�?             5@                     	          ����?���y4F�?             3@                      	          ����?�q�q�?             "@                                 �o@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                      	          ����?ףp=
�?             $@        ������������������������       �                     @                                  pc@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                +                    �?�{���l�?g            �c@       !       (                   @[@��V9��?\            �a@        "       '                    �?ףp=
�?             $@       #       $                    �?؇���X�?             @       ������������������������       �                     @        %       &                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        )       *       	             @��"pK�?V            ``@       ������������������������       �        U            @`@        ������������������������       �                     �?        ,       1                    �?      �?             0@       -       .                   �g@�<ݚ�?             "@       ������������������������       �                     @        /       0                   �h@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        3       :                    �N@���Q��?/            @P@        4       5       
             �?      �?             8@        ������������������������       �                     *@        6       7                   �d@"pc�
�?	             &@       ������������������������       �                      @        8       9                   �e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ;       N                    �?���� �?            �D@       <       =                    �?4�2%ޑ�?            �A@        ������������������������       �        	             (@        >       ?                   `[@�LQ�1	�?             7@        ������������������������       �                     @        @       E                   `a@      �?             4@        A       D                    @O@ףp=
�?             $@        B       C       	          @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        F       M                   `c@���Q��?             $@       G       L                     R@      �?              @       H       K                   �p@؇���X�?             @        I       J                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        O       P       	          ���ٿ      �?             @        ������������������������       �                     �?        Q       R                     P@���Q��?             @        ������������������������       �                      @        S       T                   `c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        V       i       
             �?�ɞ`s�?*            �N@       W       Z                    �G@؇���X�?!            �H@        X       Y                   `e@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        [       ^                    �?t��ճC�?             F@        \       ]       	             �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        _       h                    �?�(\����?             D@        `       g                   P`@��S�ۿ?             .@        a       b       
             �?r�q��?             @        ������������������������       �                      @        c       d                   Xq@      �?             @        ������������������������       �                      @        e       f                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     9@        ������������������������       �        	             (@        k       �                    �G@����&�?           Py@        l       s                   i@�,�٧��?2            �S@        m       r       	          ����?`Jj��?             ?@        n       o                    �?؇���X�?             ,@        ������������������������       �                     @        p       q                   �^@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     1@        t       �                   �c@�q�q��?             H@       u       �       
             �?�\��N��?             C@       v       {                    �F@      �?             4@       w       x                    �?@4և���?
             ,@       ������������������������       �                     (@        y       z                   pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        |       }                   �m@�q�q�?             @        ������������������������       �                     �?        ~                           �?z�G�z�?             @        ������������������������       �                      @        �       �                   p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@r�q��?
             2@       ������������������������       �                     .@        ������������������������       �                     @        �       �                    f@ףp=
�?             $@       ������������������������       �                     @        �       �       
             �?r�q��?             @        ������������������������       �                     @        �       �                   �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   P`@��J�n�?�            `t@       �       �                    �?��a�Y�?�            �i@        �       �                   �a@�'݊U�?,            �P@       �       �                   0a@�D��?            �H@        ������������������������       �                     5@        �       �                   �h@���>4��?             <@        ������������������������       �                     @        �       �                    \@      �?             8@        �       �                   �Y@�����H�?             "@        �       �                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?��S���?             .@       �       �       
             �?���|���?             &@        ������������������������       �                      @        �       �       	             �?�<ݚ�?             "@        �       �       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        �       �       	          ����?��g=��?Y            @a@        �       �                    �?�����?!            �H@        �       �                   `^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �]@�㙢�c�?             G@       �       �                   �l@�<ݚ�?             B@       �       �                   �i@��Q��?             4@       �       �                   @b@؇���X�?
             ,@       ������������������������       �                     &@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �O@      �?
             0@       ������������������������       �                     *@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                   �h@X;��?8            @V@        ������������������������       �                     ;@        �       �                    �R@Hn�.P��?%             O@       �       �                   @i@�]0��<�?$            �N@        ������������������������       �                     �?        �       �                   0p@ �.�?Ƞ?#             N@        ������������������������       �                     =@        �       �                    �J@�g�y��?             ?@        �       �       	             @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?        �       �                    �K@z��`p��?Q            @^@        �       �       	          ����?v ��?            �E@        �       �       
             �?���!pc�?             6@        �       �                   Pb@r�q��?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          `ffֿ      �?	             0@        ������������������������       �                     �?        ������������������������       �                     .@        �       �                   ``@��s����?             5@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?             0@        ������������������������       �                      @        ������������������������       �        
             ,@        �       �       
             �?����?4            �S@       �       �       	          ����?ףp=
�?!             I@        �       �                    �?�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?������?            �D@       �       �                    a@ 	��p�?             =@        ������������������������       �        	             ,@        �       �                   �v@�r����?             .@       �       �                    �M@$�q-�?
             *@        �       �                   �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   �]@      �?             <@        �       �                    [@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    _@��Q��?             4@        ������������������������       �                     @        �       �                    �?      �?             ,@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ��� @�q�q�?             "@       �       �                   �e@      �?              @       �       �                   �b@؇���X�?             @        ������������������������       �                     @        �       �                    @M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�   Np	�?���Gw{�?%P�[:�?�_]H���?.�jL��?IT�n��?
��|7�?J��8D�?!Y�B�?��Moz��?UUUUUU�?UUUUUU�?333333�?ffffff�?۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?                      �?              �?      �?                      �?��{a�?a���{�?�m۶m��?�$I�$I�?6��P^C�?(������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�-4`I/�?Kz���?�D�)͋�?t�n���?�������?�������?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        {k�4w��?qBJ�eD?      �?                      �?      �?      �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        333333�?�������?      �?      �?              �?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?                      �?jW�v%j�?,Q��+�?�������?�A�A�?      �?        Nozӛ��?d!Y�B�?              �?      �?      �?�������?�������?      �?      �?      �?                      �?      �?        333333�?�������?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        &C��6��?mާ�d�?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?t�E]t�?�E]t��?      �?      �?              �?      �?        �������?333333�?�?�������?UUUUUU�?�������?              �?      �?      �?              �?      �?      �?              �?      �?                      �?              �?      �?        t��:W�?���M1j�?:�g *�?�&��jq�?�B!��?���{��?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?y�5���?�5��P�?      �?      �?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?      �?                      �?�������?�������?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?        �%�6��?��A2���?<��;�?�;���?��[���?����??4և���?������?              �?n۶m۶�?I�$I�$�?      �?              �?      �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?�?�������?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?��v`��?�(�3J��?����X�?^N��)x�?UUUUUU�?UUUUUU�?      �?                      �?d!Y�B�?�7��Mo�?�q�q�?9��8���?ffffff�?�������?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�E(B�?�u�{���?              �?�c�1ƨ?t�9�s�?;ڼOqɠ?\2�h��?      �?        �?wwwwww�?              �?�B!��?��{���?F]t�E�?]t�E�?              �?      �?                      �?      �?        ��ˠ�?�x?r���?qG�w��?G�w��?F]t�E�?t�E]t�?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?      �?              �?      �?        �a�a�?z��y���?�������?333333�?      �?                      �?      �?      �?      �?                      �?��-��-�?H�4H�4�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?������?p>�cp�?�{a���?������?              �?�?�������?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?              �?      �?      �?      �?      �?      �?                      �?�������?ffffff�?      �?              �?      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�R�[hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKӅ�h��B�4         R       	          ����?6������?�           ��@                     
             �?��_���?�             w@                                  ph@�4�M�f�?@            �Y@        ������������������������       �                     D@                      	          ����?V��z4�?%             O@                                 �c@X�EQ]N�?            �E@                                 �`@      �?             @@       ������������������������       �        
             ,@        	                           �?�X�<ݺ?	             2@       
                           �?$�q-�?             *@                                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @                                  `]@���|���?             &@        ������������������������       �                     @                                  0e@z�G�z�?             @        ������������������������       �                     @                                  �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?�d�����?             3@        ������������������������       �                     @                                  �d@�q�q�?	             (@                     	          833�?      �?              @        ������������������������       �                      @                      
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                !       	             �(��R%��?�            �p@        ������������������������       �                      @        "       9                    @��U�=��?�            �p@       #       &                   `Q@ 7���B�?z            �g@        $       %                    `Q@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        '       *                    �?P�p�_�?u            `f@        (       )                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        +       ,                    �?��Bs�?q            �e@        ������������������������       �        (             L@        -       8                   �t@ ���J��?I            @]@       .       /                   0n@ _�@�Y�?H             ]@       ������������������������       �        ,            @R@        0       7                    �? �#�Ѵ�?            �E@       1       2                   �n@�}�+r��?             C@        ������������������������       �                     �?        3       4       	            �?�?�|�?            �B@       ������������������������       �                     A@        5       6                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        :       ?                   @E@��H�}�?0            �R@        ;       >       	          ����?8�Z$���?	             *@        <       =                   �]@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        @       I                    �?r֛w���?'             O@       A       F                   pi@�:�^���?            �F@        B       E                   @h@z�G�z�?             $@       C       D                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        G       H                   �e@ >�֕�?            �A@       ������������������������       �                    �@@        ������������������������       �                      @        J       Q                   �p@�t����?             1@       K       P                   �c@����X�?             @        L       M                    �H@�q�q�?             @        ������������������������       �                     �?        N       O       	          @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        S       t                   f@xƅd�?�            �v@        T       q                    �Q@�KM�]�?B            �\@       U       X                    �?h�)S;�??            �[@        V       W       	             @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        Y       b       
             �?88��M�?<            �Z@        Z       [                   �]@�S����?
             3@        ������������������������       �                     @        \       _                    �?      �?             (@       ]       ^                   �U@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        `       a                   @_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        c       d                    �?���7�?2             V@        ������������������������       �                     ;@        e       h                    @��GEI_�?$            �N@        f       g                   �e@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        i       n                    c@ �q�q�?             H@       j       k                   p`@����?�?            �F@       ������������������������       �                    �B@        l       m                    @M@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        o       p                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        r       s                    @R@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        u       �                   �a@�����?�            �o@       v       �       	          pff�?>a�����?f             c@        w       x                    @j���� �?             A@        ������������������������       �                     @        y       z       	          `ff�?������?             ;@        ������������������������       �                     @        {       �                    �?8����?             7@        |                           �?      �?             @       }       ~                    �M@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?������?             1@       �       �                   �`@����X�?             ,@       �       �                    �G@�θ�?
             *@        ������������������������       �                     @        �       �                    �?�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �_@��|Io��?L            �]@        �       �                   �_@@�0�!��?             A@       �       �                   �\@���!pc�?             6@        ������������������������       �                      @        �       �                    �?z�G�z�?             4@        ������������������������       �                     �?        �       �       	             @�S����?
             3@       ������������������������       �                     ,@        �       �       	          ���@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        �       �       
             �?Pq�����?8            @U@       �       �                    �?��Y��]�?6            �T@        �       �                    �?���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        3            @S@        �       �                   pq@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	             @���*��?:            �X@       �       �                    @A@*-ڋ�p�?,            @S@        ������������������������       �                     @        �       �                   s@z�7�Z�?*            @R@       �       �                   pd@�n_Y�K�?%            @P@       �       �       	          ����?p�v>��?            �G@        �       �                    �?�q�q�?             (@       �       �                   �b@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �^@�q�q�?             @        ������������������������       �                     �?        �       �       	          ����?z�G�z�?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?z�G�z�?            �A@        ������������������������       �                     0@        �       �                    �?p�ݯ��?             3@       �       �                    d@      �?
             ,@       �       �                    �?�q�q�?	             (@       �       �       	          `ff�?�q�q�?             @        ������������������������       �                     �?        �       �                    @z�G�z�?             @        ������������������������       �                      @        �       �                     M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    \@b�2�tk�?             2@        ������������������������       �                     @        �       �                   �o@      �?	             ,@       �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @F@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?              @       ������������������������       �                     @        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    [@��2(&�?             6@        ������������������������       �                      @        �       �                   �f@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  ��X�5�?��S�$e�?zӛ����?Y�B��?�������?





�?              �?�s�9��?2�c�1�?qG�wĽ?w�qG�?      �?      �?              �?�q�q�?��8��8�?;�;��?�؉�؉�?      �?      �?      �?                      �?              �?              �?F]t�E�?]t�E]�?              �?�������?�������?      �?              �?      �?      �?                      �?Cy�5��?y�5���?      �?        �������?�������?      �?      �?      �?        UUUUUU�?�������?      �?                      �?      �?        ����N��?,�T�R�?              �?�>���?|��|�?	�%����?h/�����?ffffff�?333333�?      �?                      �?B�D�H�?�7Ck��?�������?UUUUUU�?      �?                      �?s��3�q�?�������?      �?        ��-��-�?�A�A�?#,�4�r�?�{a���?      �?        �/����?�}A_Ч?�5��P�?(�����?              �?*�Y7�"�?к����?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?{�G�z�?
ףp=
�?;�;��?;�;��?�������?333333�?      �?                      �?              �?���{��?�B!��?}�'}�'�?l�l��?�������?�������?�q�q�?�q�q�?      �?                      �?              �?��+��+�?�A�A�?      �?                      �?�������?�������?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?�ݮ��?@�H�{�?(�����?�k(���?� O	�?b�־a�?UUUUUU�?UUUUUU�?      �?                      �?����f��?+J�#��?^Cy�5�?(������?              �?      �?      �?�q�q�?�q�q�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?�.�袋�?              �?;ڼOqɰ?�d����?;�;��?;�;��?              �?      �?        UUUUUU�?�������?l�l��?��I��I�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?�,˲,��?�i��i��?�?�������?ZZZZZZ�?�������?      �?        {	�%���?B{	�%��?              �?8��Moz�?d!Y�B�?      �?      �?�������?333333�?      �?                      �?      �?        �?xxxxxx�?�$I�$I�?�m۶m��?�؉�؉�?ى�؉��?              �?333333�?ffffff�?      �?                      �?      �?                      �?:�:��?��O��O�?�������?ZZZZZZ�?t�E]t�?F]t�E�?      �?        �������?�������?      �?        ^Cy�5�?(������?              �?333333�?�������?      �?                      �?              �?�?~~~~~~�?������?8��18�?�������?333333�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�@�_)�?�~�@��??!��O��?��cj`��?              �?�I�&M��?�lٲe��?;�;��?ى�؉��?ڨ�l�w�?L� &W�?�������?�������?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?�������?      �?        ^Cy�5�?Cy�5��?      �?      �?�������?�������?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?      �?                      �?      �?              �?        9��8���?�8��8��?              �?      �?      �?�������?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?t�E]t�?��.���?      �?        �������?ffffff�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�v}hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKͅ�h��B@3         x                    �?U�ք�?�           ��@                                  �?~e�.y�?
            z@                                  �Q@d�.����?K            @^@        ������������������������       �                     @                      
             �?t��%�?H            �\@                                   �?��R[s�?            �A@                                 `X@     ��?             @@        ������������������������       �                      @        	       
                    @�r����?             >@       ������������������������       �                     7@                                  �a@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                  @c@�(\����?4             T@       ������������������������       �        0             R@                                   @      �?              @       ������������������������       �                     @        ������������������������       �                      @               #                   �_@�?ȇ�p�?�            pr@                                   �?j�'�=z�?)            �P@                     
             �?�e����?            �C@                     	          `ff�?�>4և��?             <@        ������������������������       �                     (@                                  `_@     ��?	             0@       ������������������������       �                     @                                  @`@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             &@                       
             �? 7���B�?             ;@       ������������������������       �        
             0@        !       "                    @I@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        $       /                    �?P�����?�            �l@        %       &                    �I@����"�?             =@        ������������������������       �                     $@        '       .                   �p@D�n�3�?
             3@       (       )                   `Q@d}h���?             ,@        ������������������������       �                     �?        *       +                   �j@8�Z$���?             *@        ������������������������       �                     @        ,       -                   �a@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        0       9                    P@��H.�!�?�             i@        1       4                    \@ףp=
�?             4@        2       3       	          �����      �?             @        ������������������������       �                     �?        ������������������������       �                     @        5       6                     O@      �?             0@       ������������������������       �                     ,@        7       8                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        :       e                   xp@<����E�?w            �f@       ;       \       	          ����?:	��ʵ�?Y            �`@       <       E                   �[@X�
����?K             ]@        =       >                   Pi@      �?             8@        ������������������������       �                     @        ?       B                   �b@���y4F�?	             3@       @       A                    @D@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        C       D                   �c@      �?              @        ������������������������       �                     @        ������������������������       �                     @        F       G                   �^@���.�6�??             W@        ������������������������       �                     ;@        H       U                    �?���Ls�?+            @P@       I       L                    @L@@4և���?#             L@       J       K                   pf@�Ń��̧?             E@       ������������������������       �                    �D@        ������������������������       �                     �?        M       T                    @M@d}h���?             ,@       N       S                    �?�q�q�?             "@       O       R                    �?���Q��?             @       P       Q                    _@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        V       [                   p@�<ݚ�?             "@       W       X                     J@      �?              @       ������������������������       �                     @        Y       Z                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ]       ^                    �E@�\��N��?             3@        ������������������������       �                     @        _       `                    `@���Q��?             .@        ������������������������       �                     @        a       b                   �`@�q�q�?             "@        ������������������������       �                     @        c       d       
             �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        f       o       
             �?k��9�?            �F@        g       l                     J@؇���X�?
             ,@       h       i       	          @33�?�8��8��?             (@       ������������������������       �                     $@        j       k                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        m       n       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        p       q                    �?��a�n`�?             ?@       ������������������������       �                     6@        r       s                    �C@�<ݚ�?             "@        ������������������������       �                     �?        t       w                     @      �?              @        u       v                    d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        y       �                    �?��Dl<�?�            �s@        z              
             �?�X����?             6@       {       |                    �K@��
ц��?	             *@        ������������������������       �                     @        }       ~                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                   �b@��(�2Y�?�            �r@       �       �                   �U@���D�k�?�            �p@        ������������������������       �                     @        �       �                    _@p-*<�(�?�            pp@       �       �                   8s@F|/ߨ�?`            @d@       �       �                    `@�k.s�׌?S            �a@        �       �                   �o@P�Lt�<�?             C@       ������������������������       �                    �@@        �       �                    �O@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        =            �Y@        �       �       
             �?؇���X�?             5@        �       �                    �R@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �t@�KM�]�?             3@        �       �                   �`@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        �       �       
             �?L��/�/�?C            @Y@       �       �                    \@������?;            @V@        �       �                   ph@d}h���?             ,@        ������������������������       �                     @        �       �                   �b@�q�q�?             "@       �       �                     I@և���X�?             @        ������������������������       �                      @        �       �       	             �?z�G�z�?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �b@Х-��ٹ?0            �R@       �       �       	          ����?@��8��?!             H@        ������������������������       �                     6@        �       �                    �? ��WV�?             :@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        �       �                    c@�����H�?             ;@        �       �                   �`@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    @���N8�?             5@        �       �                     P@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             0@        �       �                    �?�q�q�?             (@        ������������������������       �                     �?        �       �                    �?���!pc�?             &@        ������������������������       �                     @        �       �                   �Y@      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��S���?             >@        �       �       
             �?      �?             (@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                     M@�E��ӭ�?
             2@       �       �                   c@�n_Y�K�?             *@        ������������������������       �                     @        �       �                    �?z�G�z�?             $@       �       �                    @K@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �E@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ᓔ��?�5�;��?��؉���?��N��N�?j�V���?Y�����?              �?�(�j��?�q�.�|�?X|�W|��?PuPu�?      �?      �?              �?�������?�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?              �?333333�?�������?      �?              �?      �?      �?                      �?��;M��?{>�e���?|��|�?�|���?�A�A�?�-��-��?�m۶m��?�$I�$I�?              �?      �?      �?              �?r�q��?�q�q�?      �?                      �?      �?        h/�����?	�%����?              �?F]t�E�?]t�E�?      �?                      �?(�nY���?��"M�?�i��F�?	�=����?              �?l(�����?(������?I�$I�$�?۶m۶m�?              �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?=
ףp=�?��Q���?�������?�������?      �?      �?      �?                      �?      �?      �?              �?      �?      �?              �?      �?        �[�[�??�>��?��O��O�?l�l��?	�=����?���=��?      �?      �?              �?6��P^C�?(������?]t�E�?F]t�E�?              �?      �?              �?      �?              �?      �?        ���7���?Y�B��?      �?        �����?z�z��?n۶m۶�?�$I�$I�?��<��<�?�a�a�?      �?                      �?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?y�5���?�5��P�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �'}�'}�?[�[��?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?      �?                      �?�c�1��?�s�9��?      �?        �q�q�?9��8���?      �?              �?      �?      �?      �?      �?                      �?              �?M0��>��?�sHM0��?�E]t��?]t�E]�?�؉�؉�?�;�;�?      �?              �?      �?      �?                      �?      �?        *�Y7�"�?�����?�RKE,�?�՝VwZ�?      �?        [�t8�~�?5f�.��?�����H�?�Hx�5�?t�n��}?"����?(�����?���k(�?              �?�������?�������?              �?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?        (�����?�k(���?      �?      �?      �?                      �?              �?[�߈�?��<�]?�?B�P�"�?ؽ�u�{�?۶m۶m�?I�$I�$�?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?      �?      �?                      �?              �?              �?O贁N�?K~��K�?UUUUUU�?UUUUUU�?              �?;�;��?O��N���?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?        �a�a�?��y��y�?�������?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?F]t�E�?t�E]t�?      �?              �?      �?      �?      �?      �?                      �?              �?�������?�?      �?      �?      �?      �?      �?                      �?      �?        r�q��?�q�q�?ى�؉��?;�;��?      �?        �������?�������?�$I�$I�?۶m۶m�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg}�XhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK녔h��B�:         �                    �?0����?�           ��@              ?       
             �?�ua��?           @{@                      	          ����?n2�`���?b            `c@                                   @�C��2(�?            �K@                                   @E@�q�q�?             .@                                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        	                           �?"pc�
�?	             &@       
                          �c@ףp=
�?             $@       ������������������������       �                     @                                  �`@      �?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     D@                                   �?Fx$(�?D             Y@                                   @      �?             4@                                 `X@      �?             0@        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     @               >                   �t@���Q8�?5             T@              1                   �`@      �?3             S@              (                   Pl@8�$�>�?            �E@                                  �?      �?             8@                                  �?����X�?
             ,@        ������������������������       �                     @        ������������������������       �                     $@                '                    �?z�G�z�?             $@       !       $       
             �?���Q��?             @        "       #       	             @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        %       &                   �h@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        )       .                    `@�S����?             3@       *       -                   �]@      �?
             0@        +       ,                    �D@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        /       0                   �q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        2       9                   c@<���D�?            �@@       3       4                   `c@���7�?             6@       ������������������������       �                     ,@        5       8                    @      �?              @        6       7       	          833�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        :       =                   �o@���!pc�?             &@        ;       <       	          ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        @       I                    �?��L��?�            �q@        A       H       	          ����?P�Lt�<�?0             S@       B       G                     Q@���#�İ?$            �M@       C       D                   �b@ _�@�Y�?#             M@       ������������������������       �                     J@        E       F                     @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        J       ]                   @E@�0]�I�?�            �i@        K       V                    @��+7��?             7@        L       Q                    �?      �?              @        M       N                    �?      �?             @        ������������������������       �                     �?        O       P                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        R       U                    �?      �?             @       S       T                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        W       X                   `[@�r����?
             .@        ������������������������       �                     �?        Y       \                    [@@4և���?	             ,@        Z       [                   �X@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ^       q                   0n@|)����?u            �f@       _       `                   �c@���7�?I            �[@       ������������������������       �        )            �M@        a       b                    �?`�H�/��?             �I@        ������������������������       �                     �?        c       n                    �L@HP�s��?             I@       d       e                    @=QcG��?            �G@       ������������������������       �                    �A@        f       g                   �g@      �?             (@        ������������������������       �                     �?        h       m                   @b@"pc�
�?             &@       i       j       	             �?ףp=
�?             $@       ������������������������       �                      @        k       l                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        o       p                    a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        r       �                    �?�ӭ�a��?,             R@       s       t                    �?�����?$            �O@        ������������������������       �                     �?        u       �       	             �?6uH���?#             O@       v       �       	          ����? 	��p�?              M@       w       �       	            �?�:�]��?            �I@       x                          �c@      �?             H@       y       z                    �?ȵHPS!�?             :@        ������������������������       �                     (@        {       ~                    @d}h���?             ,@        |       }                    @E@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     6@        �       �                    q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @K@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @X�<ݚ�?             "@       �       �                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@�q�� �?�            �r@       �       �                   P`@�A����?�            @q@       �       �       
             �?�qM�R��?~             i@       �       �       	          ����?��?}�?s             g@        �       �       	          hff�?f>�cQ�?'            �N@        ������������������������       �                     3@        �       �                    �?d}h���?             E@        ������������������������       �                     @        �       �                    @8�Z$���?            �C@        �       �                   �]@�q�q�?             "@       ������������������������       �                     @        �       �                   p`@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?ףp=
�?             >@        �       �                    @M@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �K@ ��WV�?             :@       ������������������������       �        
             1@        �       �                   �e@�����H�?             "@       ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �R@�â��,�?L             _@       �       �       	          ���@�-.�1a�?K            �^@       �       �                   �\@�����?>            @Y@        �       �                   `_@ףp=
�?             $@       ������������������������       �                      @        �       �                   �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        7            �V@        �       �                   �_@���7�?             6@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     �?        �       �                   �^@      �?             0@       �       �                     @�θ�?             *@        ������������������������       �                      @        �       �                   �`@�C��2(�?             &@       �       �                    �?r�q��?             @       �       �                     P@z�G�z�?             @       �       �       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @z�G�z�?1            �R@        �       �                   �o@���Q��?             $@        �       �       	             �?z�G�z�?             @        ������������������������       �                     @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?�z����?)            @P@       �       �                   �m@�C��2(�?#            �K@       �       �                   pa@д>��C�?             =@        ������������������������       �                     "@        �       �                   �m@      �?             4@       �       �                   `b@r�q��?             2@       �       �       	             �?�8��8��?
             (@        �       �                   �`@z�G�z�?             @        �       �                     L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     :@        �       �                   @b@���Q��?             $@       �       �                   @`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @���|���?             6@        ������������������������       �                     "@        �       �                   �d@�n_Y�K�?	             *@       �       �       
             �?z�G�z�?             $@        �       �                   pm@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�B�  ���^L�?���Y�?`�~�6�??Y����?��=��?�qa�?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?F]t�E�?/�袋.�?�������?�������?              �?      �?      �?      �?      �?      �?                      �?              �?      �?                      �?R���Q�?ףp=
��?      �?      �?      �?      �?              �?      �?                      �?ffffff�?�������?      �?      �?�5eMYS�?6eMYS��?      �?      �?�$I�$I�?�m۶m��?      �?                      �?�������?�������?333333�?�������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        ^Cy�5�?(������?      �?      �?UUUUUU�?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?|���?|���?F]t�E�?�.�袋�?              �?      �?      �?      �?      �?              �?      �?                      �?t�E]t�?F]t�E�?      �?      �?      �?                      �?              �?      �?        ����?�\���?���k(�?(�����?��N��?'u_[�?#,�4�r�?�{a���?      �?        �������?UUUUUU�?      �?                      �?              �?      �?        ٚ��I��?���Iٚ�?Y�B��?zӛ����?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�?�������?      �?        �$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?              �?      �?                      �?��/��/�?h�h��?�.�袋�?F]t�E�?      �?        �������?�?              �?q=
ףp�?{�G�z�?x6�;��?AL� &W�?      �?              �?      �?              �?/�袋.�?F]t�E�?�������?�������?      �?              �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�8��8��?=��<���?�a�a�?              �?k���Zk�?��RJ)��?������?�{a���?}}}}}}�?�?      �?      �?��N��N�?�؉�؉�?      �?        I�$I�$�?۶m۶m�?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?�q�q�?r�q��?�������?�������?      �?                      �?              �?�=l}0�?�� ���?�Mozӛ�?C���,�?���@��?�n�Wc"�?�	A����?��ׄ���?�u�y���?��!XG�?              �?۶m۶m�?I�$I�$�?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?�������?      �?      �?      �?                      �?;�;��?O��N���?              �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?�c�1Ƙ?:�s�9�?�h
���?{����z�?��be�F�?�tj��?�������?�������?              �?      �?      �?      �?                      �?              �?F]t�E�?�.�袋�?      �?      �?      �?                      �?              �?      �?              �?      �?�؉�؉�?ى�؉��?      �?        F]t�E�?]t�E�?UUUUUU�?�������?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?      �?        �������?�������?�������?333333�?�������?�������?      �?              �?      �?              �?      �?                      �?�Z��Z��?[��Z���?F]t�E�?]t�E�?|a���?a���{�?              �?      �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?333333�?�������?�������?�������?      �?                      �?      �?        ]t�E]�?F]t�E�?      �?        ى�؉��?;�;��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	�tlhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�-         X                    @�+	G�?�           ��@               5       
             �?bPD΂_�?�            �u@                                  �a@�zv�X�?T            �`@                                   �?     ��?*             P@                                 p`@�������?             A@                                 `X@8�A�0��?             6@        ������������������������       �                      @               	                   �X@X�Cc�?             ,@        ������������������������       �                      @        
                           �?�q�q�?
             (@        ������������������������       �                      @                                   `@      �?             $@                                  �?      �?              @                                 `]@      �?             @        ������������������������       �                      @                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@                                  P`@(;L]n�?             >@                      	             �?�����H�?             "@       ������������������������       �                     @                                  �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@               *                   �n@<��¤�?*             Q@              #                   �\@���!pc�?             F@               "                    �?      �?              @               !       	          ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        $       '       	          `ff@r�q��?             B@       %       &                   Pg@     ��?             @@        ������������������������       �                     @        ������������������������       �                     =@        (       )                    W@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        +       0                    �?      �?             8@        ,       /                    �?؇���X�?             @        -       .                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        1       4       	             �?@�0�!��?	             1@        2       3                    ^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        6       7                   �O@��$xtW�?�            �j@        ������������������������       �                     @        8       A                    �?@�S�1�?�             j@        9       >                   �c@�θ�?
             *@       :       ;                    �P@�����H�?             "@       ������������������������       �                     @        <       =                   �a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       @                    @M@      �?             @       ������������������������       �                      @        ������������������������       �                      @        B       W                   �g@`�(c�?v            �h@       C       D                   �k@`�E���?u            @h@        ������������������������       �        1            �R@        E       T                    _@0x�!���?D            �]@        F       Q                    @L@��p\�?            �D@       G       H                    �?P�Lt�<�?             C@        ������������������������       �                     &@        I       P                    �? 7���B�?             ;@       J       O                    c@���7�?             6@        K       N                   �\@z�G�z�?             @        L       M                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                     @        R       S                    @O@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        U       V       	          833@�(�Tw�?)            �S@       ������������������������       �        (            @S@        ������������������������       �                     �?        ������������������������       �                      @        Y       p                   @E@��4:���?�            Px@        Z       o                   �`@\�t��Y�??            �Y@       [       l                   P`@� ���?0            @S@       \       c       
             �?(N:!���?,            �Q@       ]       ^                    @O@h�����?$             L@       ������������������������       �                     F@        _       b                    �O@r�q��?	             (@        `       a                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        d       g                    �J@և���X�?             ,@        e       f                   @]@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        h       k       	          ����?�z�G��?             $@        i       j                   �]@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        m       n                   �\@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     :@        q       �                    c@Pk��?�            �q@       r       �       
             �?�r����?�             l@       s       |                   �\@05D�b7�?�            �i@        t       {                   �[@�q�q�?             8@       u       v                    �?�㙢�c�?             7@       ������������������������       �        
             ,@        w       z                    �?X�<ݚ�?             "@        x       y       	             �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        }       �                   �`@�~
	�?v            �f@        ~       �                    �L@$�q-�?1            �S@              �       	          033@0�)AU��?             �L@       ������������������������       �                     K@        �       �                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @M@���N8�?             5@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?r�q��?             2@        ������������������������       �                     @        �       �                    �?      �?	             (@        �       �                    `@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   Xs@@�n���?E            �Y@       ������������������������       �        ;             V@        �       �                   �s@��S�ۿ?
             .@        ������������������������       �                     �?        ������������������������       �        	             ,@        �       �                   �`@ףp=
�?             4@        �       �                   ``@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             &@        �       �                    �?N1���?#            �N@       �       �                    �M@b�2�tk�?              K@       �       �                    @H@r٣����?            �@@       �       �                    �F@���Q��?             4@       �       �                     E@     ��?
             0@       �       �                    �B@X�<ݚ�?             "@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �e@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    �?�ՙ/�?             5@        �       �       
             �?���|���?             &@        ������������������������       �                     @        �       �                    �?      �?              @       �       �                    a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?ףp=
�?             $@        ������������������������       �                     @        �       �       	          `ff�?z�G�z�?             @        �       �                   xu@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  ��C�l�?z?+^���?tS�G�?�Y�p�?�袋.��?��.���?      �?      �?�������?�������?/�袋.�?颋.���?              �?%I�$I��?�m۶m��?      �?        �������?�������?      �?              �?      �?      �?      �?      �?      �?              �?      �?      �?              �?      �?                      �?      �?                      �?�?�������?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?KKKKKK�?iiiiii�?F]t�E�?t�E]t�?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?      �?        �������?UUUUUU�?      �?      �?              �?      �?              �?      �?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        �������?ZZZZZZ�?      �?      �?              �?      �?                      �?����?��n�?�?              �?G�<��?P���?�?ى�؉��?�؉�؉�?�q�q�?�q�q�?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?��)x9�?և���X�??��W�?����?      �?        ��~���?�5�5�?�]�ڕ��?��+Q��?���k(�?(�����?      �?        	�%����?h/�����?�.�袋�?F]t�E�?�������?�������?      �?      �?              �?      �?              �?              �?              �?        UUUUUU�?UUUUUU�?              �?      �?        p��o���?�A�A�?      �?                      �?              �?���߼��?Z�Ȑ��?��VCӽ?P ���E�?��O����?L�S�?�A�A�?|�W|�W�?�$I�$I�?�m۶m��?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?333333�?ffffff�?333333�?�������?      �?                      �?              �?�$I�$I�?۶m۶m�?              �?      �?                      �?fI9 2�?}���w��?�?�������?��߁��? ~�w �?�������?UUUUUU�?d!Y�B�?�7��Mo�?              �?�q�q�?r�q��?�������?�������?      �?                      �?              �?      �?        >)7ͣ?�o��.��?;�;��?�؉�؉�?p�}��?��Gp�?              �?UUUUUU�?UUUUUU�?      �?                      �?��y��y�?�a�a�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?              �?      �?      �?      �?      �?      �?                      �?              �?��,�?\mMw��?              �?�?�������?      �?                      �?�������?�������?9��8���?�q�q�?      �?                      �?      �?        �:ڼO�?�}�K�`�?�8��8��?9��8���?>���>�?|���?333333�?�������?      �?      �?�q�q�?r�q��?�������?�������?      �?                      �?              �?      �?              �?      �?              �?      �?              �?        �a�a�?�<��<��?]t�E]�?F]t�E�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?              �?�������?�������?      �?      �?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ޡhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK߅�h��B�7         �                    �?6������?�           ��@              c       	          ����?�C�"��?"           �{@                                 `_@n(��"�?�            v@                                   �?��
ц��?.            @P@        ������������������������       �        
             1@                                   @K@      �?$             H@               
       
             �?r�q��?             8@               	       
             �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@                      	             �?$�q-�?             *@       ������������������������       �        
             (@        ������������������������       �                     �?                      
             �?�q�q�?             8@                                 8w@�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?                                   @M@�q�q�?             @        ������������������������       �                      @                                   �N@      �?             @        ������������������������       �                      @        ������������������������       �                      @               $                    �?F��ӭ��?�             r@               !                    �?�}#���?6            �T@                                  @p�|�i�?0             S@       ������������������������       �        )             P@                                   �r@      �?             (@                                  ^@ףp=
�?             $@                      
             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        "       #       
             �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        %       :       
             �?B�黀;�?�            �i@        &       -       	          ����?ҳ�wY;�?            �I@       '       ,                    �?��S�ۿ?             >@       (       +                    �?ףp=
�?             4@        )       *                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     $@        .       9                    @O@���N8�?             5@       /       0                    �G@X�Cc�?
             ,@        ������������������������       �                     @        1       8       	          ����?X�<ݚ�?             "@       2       3                    �?�q�q�?             @        ������������������������       �                     �?        4       7                   �l@z�G�z�?             @        5       6                   `b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ;       X       	            �?T����?c            @c@       <       U                   �g@�C����?[            �a@       =       R                   xt@��*��?Y            `a@       >       E                   `\@���}��?W            �`@        ?       D                    @F@���y4F�?             3@        @       C                    �E@և���X�?             @       A       B                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        F       K                    @���U�?J            �\@       G       J                    _@@uvI��??            �X@        H       I                   �^@(;L]n�?             >@       ������������������������       �                     =@        ������������������������       �                     �?        ������������������������       �        +             Q@        L       Q                   �q@     ��?             0@       M       P                    @E@�r����?
             .@        N       O                   �e@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        S       T                    b@      �?             @        ������������������������       �                     @        ������������������������       �                     @        V       W                    d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Y       b                    �?�eP*L��?             &@       Z       a                    �O@�q�q�?             "@       [       `                    �L@և���X�?             @       \       _                    l@z�G�z�?             @        ]       ^                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        d       w                    @���?>            @V@        e       f                    U@
;&����?             G@        ������������������������       �                     "@        g       h                   `\@�Gi����?            �B@        ������������������������       �                     @        i       v       
             �?�q�q�?            �@@       j       s                   p@
;&����?             7@       k       l                   �g@      �?             (@        ������������������������       �                     �?        m       n                   �`@"pc�
�?
             &@       ������������������������       �                     @        o       p                    @I@      �?             @        ������������������������       �                     �?        q       r                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        t       u                   �z@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        x       }       
             �?X�EQ]N�?             �E@        y       |                    �?����X�?             @       z       {                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ~       �                   pc@�8��8��?             B@              �                    �? 7���B�?             ;@        �       �                   �p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        �       �                   xu@�<ݚ�?             "@       �       �                   o@      �?              @       �       �                   �]@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?v���a�?�            @r@        �       �                    �?03�Z*!�?L            �^@        �       �       	          ����?���|���?             6@        �       �                   ``@�z�G��?             $@        �       �       
             �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �`@�q�q�?             (@        �       �                   �d@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `d@0�W���??            @Y@       �       �                   �W@�*v��?=            @X@        ������������������������       �                     �?        �       �                    l@      �?<             X@       �       �                   �b@ �h�7W�?"            �J@       �       �                   @a@����?�?            �F@       ������������������������       �                    �@@        �       �                     @�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �       
             �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �l@RB)��.�?            �E@        ������������������������       �                     �?        �       �                    �?��s����?             E@       �       �                   �s@�������?             >@       �       �                     P@�J�4�?             9@       �       �                    @���y4F�?             3@        ������������������������       �                      @        �       �                    `@�t����?             1@       �       �                   �n@"pc�
�?             &@        ������������������������       �                     �?        �       �                    �?ףp=
�?             $@       �       �                     M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @^@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @I@�8��8��?             (@        �       �                   @`@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?$�q-�?r             e@       �       �                    �? �Cc}�?J             \@        �       �       	             @���Q��?             $@       �       �                   �f@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �`@�:�]��?E            �Y@       �       �                   p@`����֜?0            �Q@       ������������������������       �        "             I@        �       �                   pp@P���Q�?             4@        ������������������������       �                     �?        ������������������������       �                     3@        �       �                    @N@     ��?             @@       �       �                    �?�q�q�?             5@       �       �                   @M@��Q��?             4@        ������������������������       �                     @        �       �       	             @������?             1@       �       �                    @L@���Q��?             $@       �       �                    @      �?              @        ������������������������       �                     �?        �       �                    �I@؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �R@0�)AU��?(            �L@       ������������������������       �        '             L@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��X�5�?��S�$e�?%`%`�?�?ݵ?��?�lK���?��'i�"�?�;�;�?�؉�؉�?      �?              �?      �?UUUUUU�?UUUUUU�?F]t�E�?]t�E�?      �?                      �?�؉�؉�?;�;��?      �?                      �?�������?UUUUUU�?�q�q�?��8��8�?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �q�q�?��8��8�?Y1P�M�?4u~�!��?�k(����?^Cy�5�?      �?              �?      �?�������?�������?�������?�������?              �?      �?              �?                      �?۶m۶m�?�$I�$I�?              �?      �?        �w ~��?<��;�?�������?�������?�?�������?�������?�������?�$I�$I�?�m۶m��?              �?      �?                      �?              �?�a�a�?��y��y�?%I�$I��?�m۶m��?      �?        �q�q�?r�q��?UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?                      �?      �?                      �?      �?        25�wL�?qV~B���?T�ik���?_���?4,�T�w�?c�>ZMB�?4�τ?�?���̮?6��P^C�?(������?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?      �?        	�#����?p�}��?�Cc}h��?9/���?�������?�?      �?                      �?      �?              �?      �?�������?�?      �?      �?      �?                      �?      �?                      �?      �?      �?              �?      �?              �?      �?      �?                      �?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?�������?�������?      �?      �?              �?      �?              �?                      �?      �?                      �?7��Mmj�?e%+Y�J�?�Mozӛ�?Y�B��?              �?o0E>��?#�u�)��?              �?UUUUUU�?UUUUUU�?Y�B��?�Mozӛ�?      �?      �?              �?/�袋.�?F]t�E�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?t�E]t�?F]t�E�?              �?      �?              �?        qG�wĽ?w�qG�?�$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?h/�����?	�%����?      �?      �?      �?                      �?              �?�q�q�?9��8���?      �?      �?      �?      �?              �?      �?                      �?      �?        �4iҤI�?ٲe˖-�?!�M!�?��~Y��?]t�E]�?F]t�E�?ffffff�?333333�?�������?333333�?              �?      �?              �?        �������?�������?      �?      �?      �?                      �?              �?���g��?�&��?�i�n�'�?��Id��?      �?              �?      �?"5�x+��?��sHM0�?l�l��?��I��I�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        ���)k��?S֔5eM�?      �?        �a�a�?z��y���?�������?�������?{�G�z�?�z�G��?(������?6��P^C�?      �?        �?<<<<<<�?F]t�E�?/�袋.�?      �?        �������?�������?�������?�������?              �?      �?                      �?              �?              �?333333�?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        ;�;��?�؉�؉�?۶m۶m�?%I�$I��?�������?333333�?�������?�������?              �?      �?                      �?�?}}}}}}�?�A�A�?�������?              �?�������?ffffff�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?ffffff�?�������?      �?        �?xxxxxx�?�������?333333�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?                      �?              �?              �?p�}��?��Gp�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJQY%hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKŅ�h��B@1         p                    �?�Z���?�           ��@              A                    @~�Q7:�?           �z@              &       
             �?X�@��l�?�            �p@                                   @B@�EH,���?4            �R@        ������������������������       �                     @                                   �?�xGZ���?1            �Q@                      	          ����?H%u��?             9@                                   c@      �?             (@       	                           �?ףp=
�?             $@        
                          �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@                                    E@�L�lRT�?"            �F@        ������������������������       �                     @                                   �?������?            �D@                     	             �?���|���?             6@                                  �^@���Q��?             $@        ������������������������       �                     @                                  �b@؇���X�?             @        ������������������������       �                     @                                  p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �h@r�q��?	             (@                                  @_@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @                !                   �b@���y4F�?             3@       ������������������������       �                     $@        "       #                    �I@X�<ݚ�?             "@        ������������������������       �                     @        $       %                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        '       >                     R@��A� �?|             h@       (       =                   h@`h���?y            �g@       )       2                    @L@�tVV�?x            �g@       *       +                   @n@ I!�}�?`            �b@       ������������������������       �        ;            �U@        ,       -                    �?��v$���?%            �N@       ������������������������       �                     F@        .       1                   @c@�IєX�?
             1@        /       0                   0o@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        3       8                    �?z�G�z�?             D@        4       7                   `q@p�ݯ��?             3@       5       6                    �M@      �?             ,@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        9       :                   �_@���N8�?             5@        ������������������������       �                     &@        ;       <                   �`@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ?       @                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        B       a       	          ����?�Q����?c             d@       C       J       
             �?\�����?A            �[@        D       E                    @M@`���i��?             F@       ������������������������       �                    �B@        F       G                   Pk@؇���X�?             @       ������������������������       �                     @        H       I                   0b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        K       P                   @E@�GN�z�?(            �P@        L       O                   �_@z�G�z�?             $@       M       N                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        Q       Z                    b@      �?              L@       R       Y                   �_@ "��u�?             I@       S       V                    �F@�LQ�1	�?             7@        T       U                   pb@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        W       X                   �q@�X�<ݺ?             2@       ������������������������       �        
             1@        ������������������������       �                     �?        ������������������������       �                     ;@        [       \                   pc@�q�q�?             @        ������������������������       �                     �?        ]       ^                     E@z�G�z�?             @        ������������������������       �                      @        _       `                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        b       o                    @Q@�:pΈ��?"             I@       c       h                   �t@8��8���?!             H@       d       e                   pb@��Y��]�?            �D@       ������������������������       �                     >@        f       g                   �d@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        i       n                    @O@և���X�?             @       j       m                   �`@z�G�z�?             @        k       l                   �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        q       �       
             �?$��n�?�             s@       r       �                    �?��Fi�1�?�            0p@       s       �                    �J@��wv��?y             g@        t       �                   0a@���!pc�?,            @S@       u       �                   �_@PN��T'�?             K@        v       w                    @H@��+7��?             7@       ������������������������       �                     (@        x       {                    �I@�eP*L��?             &@        y       z                   �\@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        |       }                    @J@�q�q�?             @        ������������������������       �                     @        ~                          po@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    b@`Jj��?             ?@       ������������������������       �        
             0@        �       �       	             �?�r����?             .@        �       �                   �_@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?\X��t�?             7@       �       �       	          ����?X�<ݚ�?             2@       ������������������������       �                     "@        �       �                     H@�����H�?             "@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    c@�����H�?M             [@       �       �                    @�b�E�V�?J            �Y@        �       �                   �r@؇���X�?             5@       �       �                   `[@�KM�]�?             3@        �       �                    �?      �?              @       �       �       	             �?���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   h@0��P�?<            �T@        ������������������������       �                     <@        �       �       	          ����?h�WH��?*             K@        �       �       	          ����?����X�?
             ,@        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@        �       �                   �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ^@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   `i@�(\����?              D@        ������������������������       �                     �?        ������������������������       �                    �C@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �\@`׀�:M�?.            �R@        �       �                    �Q@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                      K@        �       �                    @�[�IJ�?!            �G@        ������������������������       �                     3@        �       �       	          ����?����X�?             <@        �       �                    �?և���X�?             ,@        ������������������������       �                     @        �       �                    �?z�G�z�?             $@       �       �                   @`@�����H�?             "@        ������������������������       �                     @        �       �                   �d@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    c@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  �H���x�?����C�?�@�Ե�?��~!V��?.�jL��?IT�n��?7�i�6�?�_,�Œ�?              �?�_�_�?�A�A�?)\���(�?���Q��?      �?      �?�������?�������?      �?      �?      �?                      �?      �?                      �?      �?        l�l��?�I��I��?      �?        ��+Q��?�v%jW��?F]t�E�?]t�E]�?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?      �?      �?      �?                      �?              �?(������?6��P^C�?              �?�q�q�?r�q��?              �?UUUUUU�?UUUUUU�?              �?      �?        b6�5��?�LF�W>�?�䣓�N�?p����?ڨ�l�w�?br1���?�|����?к���{?      �?        .�u�y�?;ڼOqɐ?      �?        �?�?�������?�������?              �?      �?              �?        �������?�������?^Cy�5�?Cy�5��?      �?      �?              �?      �?              �?        ��y��y�?�a�a�?      �?        �������?�������?              �?      �?                      �?      �?      �?      �?                      �?�������?333333�?A��)A�?߰�k��?F]t�E�?F]t�E�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �袋.��?]t�E�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?�G�z�?���Q��?��Moz��?Y�B��?333333�?�������?      �?                      �?��8��8�?�q�q�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �Q����?��Q���?�������?�������?������?8��18�?              �?F]t�E�?]t�E�?              �?      �?        �$I�$I�?۶m۶m�?�������?�������?      �?      �?      �?                      �?      �?                      �?      �?        �.��.��?J��I���?�Q:���?ʼk1���?Rm�J��?��Qm�J�?t�E]t�?F]t�E�?h/�����?&���^B�?Y�B��?zӛ����?              �?t�E]t�?]t�E�?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        �B!��?���{��?              �?�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?!Y�B�?��Moz��?�q�q�?r�q��?              �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?        �q�q�?�q�q�?��,�?�jch���?�$I�$I�?۶m۶m�?(�����?�k(���?      �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?              �?      �?        8��18�?���|�?              �?B{	�%��?��^B{	�?�$I�$I�?�m۶m��?              �?�q�q�?r�q��?�������?�������?      �?                      �?      �?      �?      �?                      �?�������?333333�?      �?                      �?�������?�������?              �?      �?        к����?��L��?�������?ffffff�?              �?      �?                      �?���
b�?m�w6�;�?      �?        �$I�$I�?�m۶m��?۶m۶m�?�$I�$I�?      �?        �������?�������?�q�q�?�q�q�?              �?�������?�������?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��fbhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK߅�h��B�7         V                    @�#i����?�           ��@               ;       
             �?,Tg�x0�?�             u@               *                    �?��۾%d�?L             ]@                                 �c@��Q���?3             T@                                 @e@�jTM��?&            �N@                                  �E@z�G�z�?$            �K@        ������������������������       �                     @                                   �R@H%u��?"             I@       	                          �r@�8��8��?!             H@       
              
             �?�nkK�?             G@                      	          033�?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                      	          `ff�?�(\����?             D@       ������������������������       �                     ?@                                  �`@�����H�?             "@                                  0b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                  @_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                      
             �?p�ݯ��?             3@        ������������������������       �                     @                                   �A@      �?             0@        ������������������������       �                     �?               )                    �?z�G�z�?             .@              $                    �?d}h���?
             ,@               #                    d@�C��2(�?             &@        !       "                   `n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        %       &                    �I@�q�q�?             @        ������������������������       �                     �?        '       (                    e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        +       ,                    �K@*O���?             B@        ������������������������       �                     *@        -       :                   �z@\X��t�?             7@       .       9                   �d@�ՙ/�?             5@       /       0                    [@��S���?             .@        ������������������������       �                      @        1       8       	          ���@�n_Y�K�?             *@       2       7                    �N@z�G�z�?             $@        3       4                    \@      �?             @        ������������������������       �                     �?        5       6       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        <       E                   `_@�L�3�?�            �k@        =       >                    ^@�q�q�?             8@       ������������������������       �                     (@        ?       @                   ``@�q�q�?             (@        ������������������������       �                      @        A       D                    �?z�G�z�?             $@        B       C                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        F       U       	          ���@�ib�=�?r            �h@       G       N                    @L@��KL�6�?o            �g@       H       M                   @[@�1���܋?W            @b@        I       J                    �F@@4և���?             ,@       ������������������������       �                     "@        K       L                   @c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        R            �`@        O       R                   �_@Du9iH��?            �E@        P       Q       	          @33�?      �?              @       ������������������������       �                     @        ������������������������       �                      @        S       T                   @t@��?^�k�?            �A@       ������������������������       �                     A@        ������������������������       �                     �?        ������������������������       �                     @        W       p                   �_@D�X%��?           �x@        X       c       
             �? (��?H            @\@       Y       Z       	          033�? Df@��?7            �T@       ������������������������       �        "            �I@        [       \                   �U@      �?             @@        ������������������������       �                     �?        ]       b                    `@�g�y��?             ?@        ^       a                    �?��S�ۿ?	             .@        _       `                    @N@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     0@        d       k       	          ����?r�q��?             >@        e       j                    �K@���Q��?             @       f       g                    �F@�q�q�?             @        ������������������������       �                     �?        h       i       	          `ffֿ      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        l       o                    �?HP�s��?             9@        m       n       	             �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             4@        q       �                   �`@���c��?�            �q@       r       �                    �?д>��C�?b             b@       s       �                    @L@F�t�K��?M            �\@       t       �                   �q@�����H�?-             R@       u       �                    @H@>a�����?             �I@        v       }       	             �?�q�q�?	             (@        w       x                   �\@�q�q�?             @        ������������������������       �                     �?        y       z                   �^@z�G�z�?             @        ������������������������       �                     @        {       |                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ~                           �G@r�q��?             @       ������������������������       �                     @        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �H@$�q-�?            �C@        �       �                   �`@z�G�z�?             @        ������������������������       �                      @        �       �                   pi@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @K@�IєX�?             A@        ������������������������       �        
             1@        �       �                   @l@�t����?
             1@       ������������������������       �                     &@        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        �       �                    �?�q�q�?              E@        ������������������������       �                     @        �       �       	             �?���"͏�?            �B@        �       �                   �Z@؇���X�?             @       ������������������������       �                     @        �       �                   Pj@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �L@ףp=
�?             >@        �       �                    ^@      �?             @        ������������������������       �                      @        �       �                   �`@      �?             @        �       �                   `Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        �       �                   �h@��a�n`�?             ?@        �       �                   �Y@���Q��?             @        �       �                   �W@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �Y@ ��WV�?             :@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        �       �       
             �?�8p/�5�?Y            �a@       �       �                    @L@ДX��?.             Q@        �       �                   �\@@-�_ .�?            �B@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             @@       ������������������������       �                     <@        �       �                   (p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �m@�חF�P�?             ?@        �       �                   Pb@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�nkK�?             7@        �       �                   �c@r�q��?             @        �       �                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        �       �       	          ����?�E��ӭ�?+             R@       �       �                    �L@Z���c��?%            �O@       �       �                    �?8��8���?             H@       �       �       	          ����?�Ra����?             F@       �       �                    ]@$G$n��?            �B@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   pf@�g�y��?             ?@       ������������������������       �                     ;@        �       �                   �f@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �N@��S���?	             .@        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                   f@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   pm@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �[@�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �d@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �t�b�9     h�h)h,K ��h.��R�(KK�KK��hb�B�  �5�;���?%e��?z��y���?�0�0�?a����?sO#,�4�?�������?333333�?.�u�y�?�y��!�?�������?�������?      �?        ���Q��?)\���(�?UUUUUU�?UUUUUU�?d!Y�B�?�Mozӛ�?UUUUUU�?�������?      �?                      �?�������?333333�?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ^Cy�5�?Cy�5��?              �?      �?      �?              �?�������?�������?I�$I�$�?۶m۶m�?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        �q�q�?�q�q�?      �?        ��Moz��?!Y�B�?�a�a�?�<��<��?�?�������?              �?;�;��?ى�؉��?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?      �?        =%�S�<�?־a��?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?����>4�?/�����?*��ԟR�?�Zk��?~������?���|?n۶m۶�?�$I�$I�?      �?        �������?�������?              �?      �?              �?        qG�w��?w�qGܱ?      �?      �?      �?                      �?_�_��?�A�A�?      �?                      �?              �?R@�O.D�?�ol���?x�!���?H���?��k���?c��7�:�?              �?      �?      �?      �?        �B!��?��{���?�?�������?�������?�������?              �?      �?                      �?              �?UUUUUU�?�������?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        {�G�z�?q=
ףp�?�������?333333�?              �?      �?                      �?�-q����?i�
���?|a���?a���{�?:��,���?1��t��?�q�q�?�q�q�?�?�������?�������?�������?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?              �?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?        ;�;��?�؉�؉�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�?�?              �?�?<<<<<<�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?        *�Y7�"�?v�)�Y7�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?      �?              �?      �?      �?      �?      �?                      �?              �?              �?�c�1Ƹ?�s�9��?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?;�;��?O��N���?�������?�������?              �?      �?                      �?�������?;��:���?ZZZZZZ�?�������?к����?S�n0E�?�������?�������?              �?      �?              �?      �?              �?      �?      �?      �?                      �?��RJ)��?�Zk����?      �?      �?              �?      �?        d!Y�B�?�Mozӛ�?UUUUUU�?�������?      �?      �?      �?                      �?              �?              �?�q�q�?r�q��?Y�eY�e�?��i��i�?�������?�������?]t�E]�?]t�E�?к����?���L�?UUUUUU�?UUUUUU�?      �?                      �?��{���?�B!��?      �?              �?      �?              �?      �?              �?              �?        �������?�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?�q�q�?9��8���?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$�phG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�-         t       
             �?"��G,�?�           ��@              +                    �?�*�@P��?            {@                                   �?�G��l��?*            �O@                                  @���|���?            �@@                                 �X@�KM�]�?             3@        ������������������������       �                     �?               
                    �?�X�<ݺ?             2@              	                   `X@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@                                    Q@����X�?
             ,@                                 �c@r�q��?	             (@                                 �n@ףp=
�?             $@       ������������������������       �                     @                                  �b@      �?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @               "                   pl@���Q��?             >@               !                   Pj@���!pc�?             &@                                  @���Q��?             @        ������������������������       �                     �?                                    �?      �?             @                     	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        #       (                   �`@���y4F�?             3@        $       '                    �?      �?             @       %       &                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        )       *                     H@��S�ۿ?	             .@        ������������������������       �                     �?        ������������������������       �                     ,@        ,       ;                   �g@\�?A�?�            0w@        -       8                   �c@���f�?L             `@       .       5                    �Q@��Y��]�?G            �^@       /       4       	             �?P����?D            �]@        0       1       	          033�? >�֕�?            �A@       ������������������������       �                     >@        2       3                   `W@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        0            �T@        6       7                   @L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        9       :                   0d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        <       U                    �?d�.����?�            @n@        =       >                   @h@z�G�z�?+            �R@        ������������������������       �                     @        ?       @                   �Q@r�q��?)             R@        ������������������������       �                      @        A       T                   0n@؇���X�?(            �Q@       B       K                   �l@      �?             D@       C       D                   �_@\-��p�?             =@        ������������������������       �        
             1@        E       J                    �?�q�q�?
             (@       F       G                   @^@      �?              @        ������������������������       �                     @        H       I                    �O@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        L       M                    m@�eP*L��?             &@        ������������������������       �                     @        N       S                    @      �?              @       O       R                    �?���Q��?             @       P       Q                    �E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     >@        V       q                    c@�^����?a            �d@       W       X                    �?�Zl�i��?]            @d@        ������������������������       �                     @        Y       `       	          ����?,_ʯ08�?\            �c@        Z       _                   �\@����X�?	             5@       [       \                   �k@���Q��?             $@        ������������������������       �                     @        ]       ^                   �r@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        a       j                   �_@@��9U��?S            @a@        b       i                   �^@V�a�� �?             =@       c       d                    @PN��T'�?             ;@        ������������������������       �                      @        e       h                   �[@�J�4�?             9@       f       g                   �k@����X�?             ,@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     &@        ������������������������       �                      @        k       l                    �?��wڝ�?B            @[@       ������������������������       �        -            �R@        m       p                   pn@��?^�k�?            �A@        n       o                   p`@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     4@        r       s                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        u       �       	             �?DE��2{�?�            �r@       v       }                    I@��ED���?�             p@        w       x                    @���y4F�?             3@        ������������������������       �                     @        y       z                    �M@      �?	             0@       ������������������������       �                     (@        {       |                   �a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ~       �                    @��n�'��?�            �m@              �                    �?x/ ��?s            �f@        ������������������������       �        )             N@        �       �                    @L@�٠n�}�?J            �^@       �       �                    @G@��s��?;            �W@       ������������������������       �                    �G@        �       �                   n@�8��8��?             H@       ������������������������       �                     >@        �       �                   �\@�<ݚ�?             2@        ������������������������       �                     @        �       �                    �?��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        �       �                    �?�+$�jP�?             ;@       �       �                     M@      �?             4@        ������������������������       �                      @        �       �                   Pc@r�q��?
             2@       �       �                    `@�t����?	             1@        �       �                   `n@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@��h!��?#            �L@        ������������������������       �                     7@        �       �                   l@��.k���?             A@        �       �                    �?d}h���?             ,@        ������������������������       �                      @        �       �                   �e@�8��8��?             (@       �       �                   �^@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �M@      �?             4@       �       �                   @c@�t����?             1@        ������������������������       �                     �?        �       �                   �q@      �?
             0@       ������������������������       �                     (@        �       �                   �_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?և���X�?             E@        �       �                    �Q@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?:ɨ��?            �@@       �       �                   @b@j���� �?             1@       �       �                    �?��
ц��?	             *@        �       �                   `T@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �Y@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             0@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  �UK���?U�)|��?��Tx*<�?���a���?1�0��?��y��y�?]t�E]�?F]t�E�?�k(���?(�����?              �?��8��8�?�q�q�?�q�q�?�q�q�?              �?      �?              �?        �$I�$I�?�m۶m��?UUUUUU�?�������?�������?�������?              �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?      �?        �������?333333�?F]t�E�?t�E]t�?�������?333333�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        (������?6��P^C�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �?�������?      �?                      �?Č��:�?hn �آ�?��=aOأ?�'�	{��?������?8��18�?'u_[�?�V'u�?�A�A�?��+��+�?              �?�������?333333�?              �?      �?                      �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?Y�����?j�V���?�������?�������?      �?        UUUUUU�?�������?      �?        �$I�$I�?۶m۶m�?      �?      �?�{a���?a����?              �?UUUUUU�?UUUUUU�?      �?      �?              �?�������?�������?      �?                      �?              �?t�E]t�?]t�E�?      �?              �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?W��1 �?ՃF��[�?�����H�?�"e����?      �?        ��J�?����6b�?�$I�$I�?�m۶m��?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?                      �?              �?�Q�g���?�ځ�v`�?a���{�?��{a�?h/�����?&���^B�?              �?{�G�z�?�z�G��?�$I�$I�?�m۶m��?      �?                      �?              �?      �?        �,�M�ɂ?N��ش�?              �?�A�A�?_�_��?�?�������?              �?      �?                      �?333333�?�������?              �?      �?        ,�Œ_,�?O贁N�?�'�	�?��=aO��?(������?6��P^C�?      �?              �?      �?              �?      �?      �?              �?      �?        ��Ϣ��?P���:Ǻ?��j��j�?�Q�Q�?      �?        Pq����?�u�y��?q�����?�X�0Ҏ�?      �?        UUUUUU�?UUUUUU�?      �?        9��8���?�q�q�?              �?�������?�?      �?                      �?/�����?B{	�%��?      �?      �?              �?�������?UUUUUU�?<<<<<<�?�?      �?      �?      �?                      �?      �?                      �?      �?        Hp�}�?p�}��?      �?        �������?�?۶m۶m�?I�$I�$�?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?              �?      �?      �?<<<<<<�?�?              �?      �?      �?      �?              �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?�q�q�?�q�q�?      �?                      �?e�M6�d�?N6�d�M�?�������?ZZZZZZ�?�؉�؉�?�;�;�?�������?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW:+LhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKӅ�h��B�4         H                   �`@�#i����?�           ��@                                   �?p�L���?�            `s@                      
             �?�X����?             F@               	                   pb@8�A�0��?             6@                                  Y@d}h���?             ,@                      	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        
                          �s@      �?              @       ������������������������       �                     @        ������������������������       �                      @                                   �?���7�?             6@                                   m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@               '       	          ����?4ԡ"���?�            �p@               &                   �c@V������?6            �R@                     
             �?�4��?/            @P@                                 �[@�KM�]�?             C@                      	          ����?     ��?             0@       ������������������������       �                     *@        ������������������������       �                     @                                  �_@���7�?             6@       ������������������������       �                     3@                      	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               !       	          ����?�q�q�?             ;@                                   @P@      �?
             0@       ������������������������       �        	             .@        ������������������������       �                     �?        "       %                   �`@���!pc�?             &@       #       $                   �[@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        (       9       	          ����?p�q��?~             h@        )       8                   �`@*
;&���?             G@       *       +                    @      �?             <@        ������������������������       �                     �?        ,       7                   @^@�<ݚ�?             ;@       -       6                    �O@�q�q�?             2@       .       5                   @o@և���X�?
             ,@       /       4                   �X@�����H�?             "@        0       3                   l@      �?             @       1       2                    \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     2@        :       E                   P`@��pBI�?_            @b@       ;       D                    �L@ ��ʻ��?Y             a@       <       C                    _@�?�|�?1            �R@        =       >                   �[@�����?             5@        ������������������������       �                     @        ?       B       	          033@�r����?             .@       @       A                    @L@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        !            �J@        ������������������������       �        (             O@        F       G                    b@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        I       �                    �?������?
           �z@       J       �                    @L@      �?�            @t@       K       x       	          033�?TWi&Ĥ�?�            `n@       L       a       
             �?�W��?�            �k@        M       R       	          ����?z�J��?            �G@        N       Q                    �?�����H�?             2@        O       P                   �c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             ,@        S       `                   �d@�c�Α�?             =@       T       [                    �?X�<ݚ�?             2@       U       Z                    @K@X�<ݚ�?             "@       V       Y                   ``@և���X�?             @       W       X                   �]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        \       ]                    @�q�q�?             "@       ������������������������       �                     @        ^       _       	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        b       i                    �D@��-��ĳ?n            �e@        c       f                    �? i���t�?#            �H@       d       e                   �S@ �#�Ѵ�?            �E@        ������������������������       �                      @        ������������������������       �                    �D@        g       h                   �\@      �?             @        ������������������������       �                     @        ������������������������       �                     @        j       o                   @[@@�n�1�?K            @_@        k       n                    @z�G�z�?             @       l       m                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        p       q                    @��d��?G             ^@       ������������������������       �        5            �W@        r       w                   ``@ ��WV�?             :@        s       t                   �_@$�q-�?	             *@       ������������������������       �                      @        u       v                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        y       �                   �_@�X����?             6@       z       {                    @C@���Q��?             $@        ������������������������       �                     @        |       }                    @H@؇���X�?             @        ������������������������       �                     @        ~       �                   �b@      �?             @              �                   pf@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �       	          ����?(Q��h�?4            @T@       �       �                     P@������?              K@       �       �                   �O@�X����?             F@        ������������������������       �                     @        �       �                   �q@      �?             D@       �       �                    �?@4և���?             <@       �       �                   Hp@�����H�?             2@       �       �                     N@      �?
             0@       ������������������������       �                     *@        �       �                   @d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?�q�q�?             (@        �       �                    �N@�q�q�?             @        ������������������������       �                     �?        �       �       	          ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?�<ݚ�?             ;@        �       �                   0b@�q�q�?
             (@        ������������������������       �                     @        �       �                   �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @P@�r����?
             .@       �       �                    �?@4և���?	             ,@        �       �                   `t@r�q��?             @        ������������������������       �                     @        �       �                   y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @��H�}�?<             Y@        �       �                   �b@r֛w���?             ?@        �       �                    �?      �?             ,@       �       �                   �o@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�IєX�?
             1@        �       �                   @`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        �       �                   @d@��X���?+            @Q@       �       �                   `\@��ɉ�?)            @P@        �       �                   @Z@���Q��?             $@        ������������������������       �                      @        �       �                   �a@      �?              @        �       �       	             �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �       	             �?�C��2(�?$            �K@        �       �                   �a@      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                    �?�q�q�?             @       �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @J@`Ql�R�?            �G@        �       �                    �?�X�<ݺ?             2@        �       �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     =@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  �5�;���?%e��?�4�M�?��,�?�E]t��?]t�E]�?/�袋.�?颋.���?۶m۶m�?I�$I�$�?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?�.�袋�?F]t�E�?      �?      �?      �?                      �?      �?        &���g¿?{����?o0E>��?�g�`�|�?�Z��Z��?�R+�R+�?(�����?�k(���?      �?      �?              �?      �?        F]t�E�?�.�袋�?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?t�E]t�?F]t�E�?�q�q�?�q�q�?      �?                      �?      �?                      �?UUUUUU�?�����*�?8��Moz�?���,d!�?      �?      �?      �?        �q�q�?9��8���?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?�q�q�?�q�q�?      �?      �?      �?      �?              �?      �?                      �?              �?      �?                      �?              �?              �?����?���Ǐ�?�?�������?к����?*�Y7�"�?�a�a�?=��<���?              �?�?�������?�$I�$I�?n۶m۶�?              �?      �?              �?                      �?              �?�������?�������?              �?      �?        �`��}�?�>����?      �?      �?��lC@��?w�M��:�?\�[��?�j��j��?}g���Q�?AL� &W�?�q�q�?�q�q�?      �?      �?              �?      �?                      �?5�rO#,�?�{a���?r�q��?�q�q�?�q�q�?r�q��?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        �f��o��?/�I���?/�����?����X�?�/����?�}A_Ч?              �?      �?              �?      �?              �?      �?        �rh��|�?����Mb�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�?      �?        O��N���?;�;��?�؉�؉�?;�;��?      �?        �������?�������?      �?                      �?      �?        ]t�E]�?�E]t��?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        x�5?,�?������?B{	�%��?{	�%���?�E]t��?]t�E]�?              �?      �?      �?n۶m۶�?�$I�$I�?�q�q�?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?        333333�?�������?              �?      �?                      �?      �?        �q�q�?9��8���?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        �?�������?�$I�$I�?n۶m۶�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        
ףp=
�?{�G�z�?���{��?�B!��?      �?      �?F]t�E�?]t�E]�?      �?                      �?      �?        �?�?UUUUUU�?UUUUUU�?              �?      �?              �?        ��v`��?�Q�g���?�����?�����?�������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?F]t�E�?]t�E�?      �?      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?W�+�ɕ?}g���Q�?�q�q�?��8��8�?      �?      �?      �?                      �?              �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJF<KdhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@/         r       
             �?�#i����?�           ��@              Q                   �b@L�~m��?           �x@                                  �?�Zl�i��?�            @t@                                  �r@�d�����?             C@              
       
             �?z�G�z�?            �A@                                   �?      �?             @        ������������������������       �                     �?               	                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �P@�חF�P�?             ?@                                  m@�r����?             >@                                  �?������?	             .@                                 �e@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                     @               N                    �R@$�q-�?�            �q@              )                    �?��d4��?�            �q@               (                    �?�q�q�?             B@                                 @[@և���X�?             <@        ������������������������       �                     @               #                   �`@�eP*L��?             6@              "                    @L@r�q��?	             (@              !                     K@�q�q�?             @                                  �a@z�G�z�?             @                                  �s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        $       %                    �?z�G�z�?             $@        ������������������������       �                     @        &       '                   p@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        *       5                    @��Ŀ�?�            �n@        +       ,                    @M@dP-���?            �G@        ������������������������       �                     5@        -       2                   �`@8�Z$���?             :@       .       1                    �M@�}�+r��?             3@        /       0       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             1@        3       4                     P@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        6       M                    �?p���?�             i@       7       L                    �?XB���?N             ]@       8       I                   @b@�kb97�?5            @S@       9       :                    @K@���(-�?1            @R@        ������������������������       �                     @@        ;       B                    `@��p\�?            �D@        <       A                   �`@"pc�
�?             &@       =       @                   �^@�q�q�?             @       >       ?                    �O@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        C       H                     L@(;L]n�?             >@        D       E                    �?ףp=
�?             $@        ������������������������       �                     @        F       G       	             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        J       K                   �h@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        ������������������������       �        9             U@        O       P                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        R       g                    �?)O���?-             R@       S       f                    �?��Q��?             D@       T       U                    K@��S���?             >@        ������������������������       �                     @        V       c                   pe@|��?���?             ;@       W       \       	          033�?���Q��?             4@       X       [                    �?z�G�z�?             $@       Y       Z       	          433�?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ]       ^                    �?���Q��?             $@        ������������������������       �                     �?        _       b                   pd@�q�q�?             "@       `       a                    @B@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        d       e                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        h       o                   0e@      �?             @@       i       j                    �L@�>4և��?             <@        ������������������������       �                     *@        k       l                    [@�q�q�?	             .@        ������������������������       �                     @        m       n       	          033�?      �?             $@        ������������������������       �                     @        ������������������������       �                     @        p       q                    @J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        s       ~                    �?4>���?�             u@        t       w                    �?���N8�?6             U@       u       v                    T@0�,���?+            �P@        ������������������������       �                      @        ������������������������       �        *            @P@        x       }                    �?�t����?             1@       y       z                    s@8�Z$���?	             *@       ������������������������       �                     "@        {       |                   �t@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               �                    @�U���?�            �o@       �       �                    @M@��C[���?c             e@       �       �                   @[@����?O            @`@        �       �                    �?և���X�?             @        ������������������������       �                     �?        �       �                   `m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    I@��Y��]�?L            �^@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �       	            �?@���a��?I            �\@       ������������������������       �        =            �W@        �       �       	          pff�?P���Q�?             4@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             2@        �       �                   ps@�	j*D�?            �C@       �       �                     R@      �?             B@       �       �                    �?     ��?             @@        �       �                     O@�eP*L��?             &@        ������������������������       �                     @        �       �       	          hff�?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     5@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?Zz�����?5            @U@       �       �                   �a@�q�q�?              H@       �       �                    X@      �?             @@        ������������������������       �                     @        �       �                    �M@XB���?             =@       ������������������������       �                     8@        �       �                    �?z�G�z�?             @       �       �                   �]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   pf@      �?             0@        ������������������������       �                     @        �       �                    �L@      �?             (@       �       �                    @F@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �J@���@��?            �B@        ������������������������       �                     &@        �       �                    @K@�	j*D�?             :@        ������������������������       �                     @        �       �                    c@��<b���?             7@       �       �                    S@ףp=
�?             4@        �       �                   �^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �5�;���?%e��?K�Z�R��?�_)P�W�?�����H�?�"e����?y�5���?Cy�5��?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��RJ)��?�Zk����?�?�������?�?wwwwww�?      �?      �?              �?      �?                      �?              �?      �?              �?        ;�;��?�؉�؉�?������?��`��?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?t�E]t�?]t�E�?�������?UUUUUU�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?              �?                      �?      �?        �������?�������?              �?�������?333333�?      �?                      �?              �?T	9?��?k�o���?W�+�ɵ?�����F�?              �?;�;��?;�;��?(�����?�5��P�?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?                      �?{�G�z�?\���(\�?�{a���?GX�i���?�cj`?�Y�	qV�?�P�B�
�?��իW��?              �?��+Q��?�]�ڕ��?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?                      �?�?�������?�������?�������?              �?�������?�������?      �?                      �?              �?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?      �?                      �?9��8���?��8��8�?ffffff�?�������?�������?�?              �?{	�%���?	�%����?�������?333333�?�������?�������?�������?333333�?      �?                      �?              �?333333�?�������?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?              �?      �?      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?��]�`��?�T�6|��?��y��y�?�a�a�?Ez�rv�?g��1��?              �?      �?        <<<<<<�?�?;�;��?;�;��?      �?              �?      �?              �?      �?              �?        ��`0�?����|>�?�wɃg�?�B���Ǽ?n�Fn�F�?�����?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?8��18�?������?      �?      �?      �?              �?      �?              �?      �?        �uI�ø�?���ρ?      �?        ffffff�?�������?      �?      �?              �?      �?              �?        vb'vb'�?;�;��?      �?      �?      �?      �?]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?      �?                      �?      �?              �?      �?      �?                      �?              �?�������?000000�?�������?�������?      �?      �?              �?GX�i���?�{a���?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?      �?      �?      �?              �?      �?                      �?к����?L�Ϻ��?              �?;�;��?vb'vb'�?      �?        ��Moz��?��,d!�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJؽ�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKׅ�h��B�5         V                    @�/�$�y�?�           ��@               ;       
             �?0�����?�            pu@               $                    �?�*;L�?N             ^@              #                   0r@rr�J��?0            �R@                                 d@.Lj���?,             Q@                     
             �?��<b���?             G@        ������������������������       �                     @                                   �?�T|n�q�?            �E@       	              	          `ff�?�'�`d�?            �@@       
                           �O@8����?             7@                                 `\@z�G�z�?             4@        ������������������������       �                     "@                                   �?���|���?	             &@                                  g@      �?              @        ������������������������       �                      @                                   @F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     $@                                   �?8�A�0��?             6@                                 pe@d}h���?
             ,@        ������������������������       �                      @                                  �`@      �?             @        ������������������������       �                     @        ������������������������       �                     @               "                    o@      �?              @              !                   �k@؇���X�?             @                                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        %       &                    \@�㙢�c�?             G@        ������������������������       �                     �?        '       2                   Pk@���V��?            �F@       (       +                    �?z�G�z�?             9@        )       *                    `@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ,       -       	          ����?ףp=
�?             4@        ������������������������       �                     $@        .       /       
             �?z�G�z�?             $@        ������������������������       �                     @        0       1                   �`@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        3       4                    @M@ףp=
�?             4@       ������������������������       �                     (@        5       6                   �`@      �?              @        ������������������������       �                     �?        7       8                   0`@؇���X�?             @       ������������������������       �                     @        9       :                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        <       U       	          ���@h�qVhԳ?�            �k@       =       D                    @L@Ц�f*�?�            �k@       >       C                    �?@�:;��?h            �f@       ?       @                   h@���1��?>            �Z@       ������������������������       �        <            �Y@        A       B                   pn@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        *            �R@        E       T                   �s@�ݜ�?            �C@       F       O       	            �?�KM�]�?             C@       G       N                    �?��S�ۿ?             >@       H       M                   �p@�����?             5@       I       J                    �Q@P���Q�?             4@       ������������������������       �                     ,@        K       L       	          ����?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        P       S                   a@      �?              @        Q       R                    �O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        W       �       	          ����?@�0�!��?�            px@        X       g                   �e@�lg����?Z             `@        Y       f                    �?(N:!���?            �A@       Z       c                   @b@���y4F�?             3@       [       b                    �?      �?             0@       \       a                    �?�<ݚ�?             "@       ]       ^       
             �?�q�q�?             @        ������������������������       �                     @        _       `       	          @33�?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        d       e       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             0@        h       �                    �?JJ����?B            �W@       i       |                   �p@��
ц��?6            �S@       j       m       
             �?��}*_��?$             K@        k       l       	          833�?�d�����?             3@       ������������������������       �        	             ,@        ������������������������       �                     @        n       {       	            �?b�h�d.�?            �A@       o       z                   �b@     ��?             @@       p       u                   �o@`Jj��?             ?@       q       r                    �? 7���B�?             ;@       ������������������������       �                     9@        s       t                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        v       w                    �?      �?             @        ������������������������       �                      @        x       y                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        }       �                    e@�q�q�?             8@       ~       �                    �?���!pc�?             6@               �                    @M@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?@�0�!��?             1@       ������������������������       �                     $@        �       �                    �I@և���X�?             @       �       �                    �?���Q��?             @       �       �                   0d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �G@      �?             0@        ������������������������       �                     �?        �       �                   �`@��S�ۿ?             .@       ������������������������       �                     $@        �       �                   `a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �R@���I���?�            `p@       �       �                   @l@(h�1W�?�            @p@       �       �                    �?0Ƭ!sĮ?T             `@        ������������������������       �                    �@@        �       �                    \@ �q�q�??             X@        �       �                    �?�q�q�?             @        �       �                   �X@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   P`@����?�?9            �V@       ������������������������       �        ,            �Q@        �       �                   �^@ףp=
�?             4@        �       �       	          033@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          033�?�IєX�?             1@        �       �                   �b@r�q��?             @        ������������������������       �                     @        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �       	          ����?HX���?M            ``@        �       �                   @_@��P���?            �D@        �       �                   �\@���Q��?             $@        ������������������������       �                      @        �       �                    @G@      �?              @       �       �                   �m@      �?             @        ������������������������       �                     �?        �       �                    b@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�חF�P�?             ?@       �       �                   �t@�q�q�?             8@       �       �                    �?؇���X�?             5@        ������������������������       �                     �?        �       �                   �`@ףp=
�?
             4@       �       �                    �N@z�G�z�?             $@       �       �                   `c@����X�?             @       �       �                    �?���Q��?             @       �       �                   hp@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                   ``@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       	             @��S�ۿ?4            �V@       �       �       	          ����? �.�?Ƞ?#             N@        �       �                     H@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �        
             0@        ������������������������       �                    �E@        �       �       	          ���@r�q��?             >@        ������������������������       �                      @        �       �                   �\@ �Cc}�?             <@        �       �                    �K@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     3@        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  L�f���?Z�L��?��Ö�j�?��xҊ*�?�������?""""""�?L�Ϻ��?Z7�"�u�?�������?------�?��Moz��?��,d!�?      �?        6eMYS��?���)k��?'�l��&�?6�d�M6�?8��Moz�?d!Y�B�?�������?�������?              �?F]t�E�?]t�E]�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?              �?颋.���?/�袋.�?I�$I�$�?۶m۶m�?      �?              �?      �?      �?                      �?      �?      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?              �?        d!Y�B�?�7��Mo�?      �?        �>�>��?[�[��?�������?�������?333333�?�������?              �?      �?        �������?�������?              �?�������?�������?              �?�$I�$I�?�m۶m��?              �?      �?        �������?�������?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?���a��?O���橤?!O	� �?�־a�?Y]����?�rS�<�v?�S�rp��?�+J�#�?      �?              �?      �?      �?                      �?      �?        \��[���?�i�i�?�k(���?(�����?�������?�?=��<���?�a�a�?ffffff�?�������?      �?        �������?UUUUUU�?              �?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?�������?ZZZZZZ�?�}A_��?}A_��?�A�A�?|�W|�W�?(������?6��P^C�?      �?      �?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?x6�;��?��
br�?�;�;�?�؉�؉�?_B{	�%�?B{	�%��?y�5���?Cy�5��?              �?      �?        ;��:���?_�_��?      �?      �?���{��?�B!��?	�%����?h/�����?      �?              �?      �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?333333�?�������?      �?                      �?�������?ZZZZZZ�?              �?۶m۶m�?�$I�$I�?333333�?�������?      �?      �?              �?      �?                      �?              �?      �?              �?      �?      �?        �?�������?              �?�������?�������?      �?                      �?���ℴ?���co�?S+�R+��?�Z��Z��?����?����?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?l�l��?��I��I�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?�?�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?J�eDP�?7Ls�U�?�����?������?�������?333333�?      �?              �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?��RJ)��?�Zk����?�������?UUUUUU�?�$I�$I�?۶m۶m�?      �?        �������?�������?�������?�������?�$I�$I�?�m۶m��?�������?333333�?      �?      �?      �?                      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�?�������?�?wwwwww�?�?�?      �?                      �?              �?UUUUUU�?�������?      �?        ۶m۶m�?%I�$I��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �t�bub�.�      hhubh)��}�(hhhhhNhKhKhG        hh%hNhJX��vhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@*         h       
             �?���
%�?�           ��@              -                    �? ��7E��?           �z@                      	          ����?�Kǔ�{�?f            `d@                                   @E@ pƵHP�?              J@                                  pe@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     F@        	       $                   �`@��_����?F            �[@       
                           \@     8�?'             P@                                   �M@����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                  �Z@�^���U�?"            �L@        ������������������������       �                     "@                                  k@r�qG�?             H@                      	          `ff@�����?             5@                                 �^@�X�<ݺ?             2@                     
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@                                  �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   @�5��?             ;@                                  @L@      �?
             4@       ������������������������       �                     (@                                  �z@      �?              @       ������������������������       �                     @        ������������������������       �                     @                #                    b@؇���X�?             @       !       "                   �n@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        %       &       	          833�?dP-���?            �G@        ������������������������       �                      @        '       ,                    �?`Ӹ����?            �F@        (       +                   P`@r�q��?             (@        )       *                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                    �@@        .       g                   �c@�iyw	
�?�            �p@       /       \                    �?���}��?�            �p@       0       3                   �Z@��5�uԾ?{            @i@        1       2                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        4       W                   �b@������?x            �h@       5       N                   �s@���|$ö?t             h@       6       =                    �?@�c��?j            �e@        7       8       	          ����?r�q��?             2@        ������������������������       �                     "@        9       :                    `@�q�q�?             "@        ������������������������       �                     @        ;       <                    _@      �?             @        ������������������������       �                     @        ������������������������       �                     @        >       M       	          ����?�#��g1�?_            �c@        ?       @                   0k@0G���ջ?"             J@       ������������������������       �                     @@        A       F                   @n@R���Q�?             4@        B       C                   @_@�q�q�?             @        ������������������������       �                     �?        D       E                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        G       L       	          ����?�IєX�?             1@        H       K                   �`@      �?              @       I       J       	          ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �        =            @Z@        O       V                    �?r�q��?
             2@       P       S                    @���!pc�?             &@        Q       R                   @[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        T       U                    �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        X       Y                    @C@�q�q�?             @        ������������������������       �                      @        Z       [                    b@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ]       d                   �`@     �?+             P@       ^       _                   �[@@�E�x�?"            �H@        ������������������������       �                     8@        `       a                   �c@`2U0*��?             9@       ������������������������       �                     7@        b       c       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        e       f                   0a@�r����?	             .@        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                      @        i       l                    �?�˱��H�?�            �r@        j       k                    T@p�qG�?=             X@        ������������������������       �                     @        ������������������������       �        <            �V@        m       z                   �O@�G�5��?�            �i@        n       o                   `]@�eP*L��?             6@        ������������������������       �                     @        p       w       	          hff�?�\��N��?             3@        q       v                    �?"pc�
�?             &@       r       s                    @ףp=
�?             $@        ������������������������       �                     @        t       u                   �]@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        x       y                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        {       �                    �?��!w�K�?v             g@       |       �                   `\@�es�q��?f            �c@        }       �                   �m@J�8���?             =@       ~       �                    �?@4և���?	             ,@              �                    @$�q-�?             *@        ������������������������       �                     @        �       �       	          ����?؇���X�?             @       �       �                    @I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    o@���Q��?             .@        ������������������������       �                     @        �       �                   �o@      �?             (@        ������������������������       �                     @        �       �                    �?      �?              @       �       �                    @N@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @L@     �?U             `@       �       �                   �g@@��8��?=             X@       �       �                   l@��K2��?;            �W@        �       �                   �b@��Y��]�?            �D@       ������������������������       �                    �C@        �       �                   0c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        !            �J@        �       �                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@     ��?             @@        �       �                   �c@�q�q�?             (@       �       �                    �L@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?ףp=
�?             4@       �       �                    q@�r����?             .@       ������������������������       �        
             *@        ������������������������       �                      @        ������������������������       �                     @        �       �                    @X�Cc�?             <@        ������������������������       �                     $@        ������������������������       �                     2@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�
  ��\���?��Q���?:�����?q����?kq�}�?�uǋ-��?;�;��?'vb'vb�?      �?      �?              �?      �?                      �?<zel���?�B�I .�?     ��?      �?�$I�$I�?�m۶m��?      �?                      �?c:��,��?:��,���?              �?UUUUUU�?UUUUUU�?=��<���?�a�a�?��8��8�?�q�q�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?h/�����?/�����?      �?      �?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?W�+�ɵ?�����F�?      �?        l�l��??�>��?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?*g��1�?����?���̮?4�τ?�?Q`ҩy�?�������?UUUUUU�?UUUUUU�?              �?      �?        ���/M�?�n-;�?�r*�?���X���?E'�卡?�M�!��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        A����?>"'wc�?�؉�؉�?vb'vb'�?              �?333333�?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�?�?      �?      �?      �?      �?              �?      �?                      �?              �?              �?UUUUUU�?�������?t�E]t�?F]t�E�?      �?      �?              �?      �?        �q�q�?9��8���?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?     ��?9/���?և���X�?              �?{�G�z�?���Q��?              �?      �?      �?      �?                      �?�?�������?      �?                      �?      �?        l����?O���!��?UUUUUU�?�������?              �?      �?        ��v`��?�%~F��?]t�E�?t�E]t�?              �?y�5���?�5��P�?/�袋.�?F]t�E�?�������?�������?      �?        �������?�������?      �?                      �?              �?      �?      �?      �?                      �?���	A�?��	A���?��9A��?9A���?�rO#,��?|a���?n۶m۶�?�$I�$I�?�؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?              �?        �������?333333�?              �?      �?      �?      �?              �?      �?      �?      �?      �?                      �?              �?     @�?      �?UUUUUU�?UUUUUU�?��Q�٨�?W�+�Ʌ?8��18�?������?      �?              �?      �?              �?      �?              �?              �?      �?      �?                      �?      �?      �?�������?�������?�������?UUUUUU�?              �?      �?                      �?�������?�������?�������?�?      �?                      �?      �?        �m۶m��?%I�$I��?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���EhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKх�h��B@4         V       	          033�?�r,��?�           ��@              #       
             �?H;N	�	�?�             x@                                  �g@�&�5y�?J             _@                                   �?`���i��?             F@                      
             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        	                          n@��Q��?.             T@        
                           �?���|���?             F@        ������������������������       �                     $@                                  �a@��.k���?             A@                      	          ����?؇���X�?	             ,@       ������������������������       �                     (@        ������������������������       �                      @                                   �J@z�G�z�?	             4@        ������������������������       �                     @                                  p`@�IєX�?             1@                                 �_@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@               "                   pq@4?,R��?             B@                                 �p@���N8�?             5@                                  �?�t����?
             1@                                   �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@                                  (q@      �?             @        ������������������������       �                      @                !                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@        $       O       	          ����?8Ӈ���?�            `p@       %       8                    @����a�?�            �n@       &       7       	          ����?`���i��?v             f@       '       4                   h@ ���l��?g            `c@       (       +                    I@���J��?e             c@        )       *                    ^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ,       /                    �?�}��L�?c            �b@        -       .                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        0       1                    �? ���?_             b@       ������������������������       �        9             U@        2       3                    �O@��v$���?&            �N@       ������������������������       �        %             N@        ������������������������       �                     �?        5       6                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        9       J                    �?�M���?(             Q@       :       ;                   �_@�����H�?             K@        ������������������������       �                     8@        <       A                   �c@z�G�z�?             >@       =       >                    �?���7�?             6@       ������������������������       �        	             0@        ?       @                   0a@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        B       C       	          `ffֿ      �?              @        ������������������������       �                      @        D       E                   �`@      �?             @        ������������������������       �                     �?        F       I                    �I@���Q��?             @        G       H                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        K       N                   �q@X�Cc�?	             ,@       L       M                   `\@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        P       Q                    �?X�<ݚ�?             2@        ������������������������       �                      @        R       S                   �U@z�G�z�?             $@        ������������������������       �                     @        T       U                    �L@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        W       �                   �b@д>��C�?�            �u@       X       q                    �?܍�l�p�?�             r@        Y       ^       
             �?d��0u��?&             N@        Z       ]                    �?      �?             $@       [       \                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        _       p                    �?�J�4�?              I@       `       o                    �?r٣����?            �@@       a       n       
             �?�LQ�1	�?             7@       b       m                    `P@����X�?             5@       c       l                    @���y4F�?             3@       d       e                   �\@���Q��?             $@        ������������������������       �                     �?        f       g                    �?�q�q�?             "@        ������������������������       �                     @        h       i                    �?      �?             @        ������������������������       �                      @        j       k                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �        	             1@        r       s                    V@ج��w�?�            �l@        ������������������������       �                     �?        t       �                   P`@T�����?�            �l@        u       v                     F@�p ��?9            �T@        ������������������������       �                     *@        w       x       
             �?�㙢�c�?2            @Q@        ������������������������       �        	             .@        y       �                    �?�<ݚ�?)             K@       z       �                    �?�d�����?             C@       {       �                   a@��<b���?             7@       |       }                    �?�t����?             1@        ������������������������       �                     �?        ~       �                   @s@      �?             0@              �                   0i@؇���X�?             ,@        �       �       
             �?�q�q�?             @       �       �                    �?z�G�z�?             @       �       �                   �^@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                     O@�q�q�?             .@       �       �                    �?�eP*L��?             &@        ������������������������       �                      @        �       �       	          ���@�q�q�?             "@       �       �                    �H@      �?              @        ������������������������       �                     �?        �       �                    `@؇���X�?             @       ������������������������       �                     @        �       �                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             0@        ������������������������       �                     �?        �       �                   �Z@��S�ۿ?             .@        �       �                   �Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             (@        �       �       	          ����?��<�Ұ?V            `b@        �       �                    `@l�b�G��?%            �L@       ������������������������       �                    �C@        �       �       	          ����?�<ݚ�?
             2@       �       �                   �l@�8��8��?             (@        �       �                   �e@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     L@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   k@�E�����?1            �V@        �       �                    �J@ qP��B�?            �E@        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     D@        ������������������������       �                    �G@        �       �                    �L@      �?&             M@       �       �                    \@P����?             C@        ������������������������       �                      @        �       �                    U@<ݚ)�?             B@        ������������������������       �                      @        �       �                    @�������?             A@       �       �                   `c@      �?             8@       �       �                   (p@���7�?             6@       ������������������������       �                     3@        �       �                   �q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   0e@���Q��?             $@        ������������������������       �                     @        �       �                   �_@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �P@z�G�z�?             4@       �       �                    a@      �?
             0@        ������������������������       �                      @        �       �                    b@      �?              @        �       �                    �?�q�q�?             @       �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  �292ȯ�?�f����?�t���L�?��|"f�?�1�c��?:�s�9�?F]t�E�?F]t�E�?�������?�������?      �?                      �?              �?ffffff�?�������?]t�E]�?F]t�E�?      �?        �������?�?�$I�$I�?۶m۶m�?              �?      �?        �������?�������?              �?�?�?      �?      �?      �?                      �?      �?        r�q��?�8��8��?��y��y�?�a�a�?�?<<<<<<�?      �?      �?              �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?                      �?�*NHɳ�?����a�?��).��?&C��6�?F]t�E�?F]t�E�?-��,�?mЦm�?______�?�?UUUUUU�?UUUUUU�?      �?                      �?�_,�Œ�?O贁N�?�������?�������?      �?                      �?x����?����?|?      �?        .�u�y�?;ڼOqɐ?      �?                      �?      �?      �?      �?                      �?      �?        �������?<<<<<<�?�q�q�?�q�q�?      �?        �������?�������?�.�袋�?F]t�E�?      �?        �������?UUUUUU�?              �?      �?              �?      �?              �?      �?      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�m۶m��?%I�$I��?�m۶m��?�$I�$I�?              �?      �?                      �?r�q��?�q�q�?      �?        �������?�������?              �?�������?333333�?      �?                      �?|a���?a���{�?)ٵ��]�?�DɮM��?�������?�?      �?      �?r�q��?�q�q�?      �?                      �?              �?{�G�z�?�z�G��?|���?>���>�?d!Y�B�?Nozӛ��?�$I�$I�?�m۶m��?(������?6��P^C�?�������?333333�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?                      �?              �?      �?              �?                      �?              �?A�V���?�%��~�?      �?        ���.�?��!:ܟ�?��+Q��?Q��+Q�?              �?d!Y�B�?�7��Mo�?              �?�q�q�?9��8���?y�5���?Cy�5��?��Moz��?��,d!�?�������?�������?      �?              �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?      �?        �?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?[��5;j�?�7�L\��?p�}��?�Gp��?              �?�q�q�?9��8���?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?      �?              �?      �?        l�l��?P��O���?�}A_З?��}A�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?�P^Cy�?Q^Cy��?              �?��8��8�?�8��8��?              �?�������?�������?      �?      �?�.�袋�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?333333�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:9)bhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�-         v                    �?T8���?�           ��@              a                    �?�yZ����?           �z@              P       	          033�?���X�K�?�            �v@              )       
             �?����j��?�            �s@                                  `]@�ހ��?:            �W@        ������������������������       �                     6@                                   �?r�q��?.             R@                                  �c@���}<S�?             7@       	       
                   �[@z�G�z�?	             $@        ������������������������       �                     �?                                   �?�����H�?             "@        ������������������������       �                     @                                   c@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@                      	          833�?f�Sc��?            �H@                     
             �?V�a�� �?             =@        ������������������������       �                     @                                    E@ȵHPS!�?             :@                                   �C@�θ�?             *@       ������������������������       �                     "@                                  �b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@               $       	          ����?���Q��?             4@                                 �_@8�Z$���?	             *@                                  �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                !                   �c@�C��2(�?             &@       ������������������������       �                      @        "       #                   �q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        %       (                     F@؇���X�?             @        &       '                   Pp@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        *       O                   �g@��X��?�             l@       +       F                   �b@���l��?�            �k@       ,       -                    �?��d5z�?�            `i@        ������������������������       �        $             K@        .       1                    X@l������?\            �b@        /       0                   �[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        2       3                    �?d�;�s��?Y            �a@        ������������������������       �                     �?        4       =                    _@���.�d�?X            �a@        5       :                    �?�J�4�?#             I@       6       7                   @^@�����?             E@       ������������������������       �                    �B@        8       9                    �C@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ;       <                    ]@      �?              @        ������������������������       �                     @        ������������������������       �                     @        >       ?                   �c@�����?5             W@        ������������������������       �                     I@        @       A                    �?�Ń��̧?             E@        ������������������������       �                     5@        B       C                   Pt@���N8�?             5@       ������������������������       �                     2@        D       E                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        G       H                    �?���y4F�?             3@        ������������������������       �                     @        I       N                   @f@������?             .@       J       K                    �?8�Z$���?             *@       ������������������������       �                     $@        L       M                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        Q       \                   �d@0,Tg��?             E@       R       W                    �?@�0�!��?             A@        S       V                    �L@���Q��?             @       T       U                   0b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        X       [       	          `ff@ܷ��?��?             =@        Y       Z                    �?z�G�z�?             .@        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     ,@        ]       ^       
             �?      �?              @        ������������������������       �                     @        _       `                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        b       c                    Z@=��T�?1            �Q@        ������������������������       �                     "@        d       i                    _@�p����?+            �N@        e       h                    @$�q-�?             :@        f       g                    @O@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     6@        j       q       
             �?����X�?            �A@        k       n                    �?���!pc�?             &@        l       m                    �P@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        o       p                    @P@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        r       u                    �?�8��8��?             8@        s       t                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     3@        w       �                   �b@�s�ۺ�?�             s@       x       �                    �?�C��2(�?�            0q@        y       �                   �a@     ��?             @@       z       {                   @[@�X����?
             6@        ������������������������       �                      @        |       }                   P`@      �?             4@        ������������������������       �                      @        ~              	          ����?�q�q�?             (@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �R@�
�3�?�            `n@       �       �                   P`@@:��JU�?�            @n@       �       �                   pl@��Μ�V�?v             h@       ������������������������       �        @             [@        �       �                   �l@@�)�n�?6            @U@        ������������������������       �                      @        �       �       
             �?��'�`�?5            �T@        ������������������������       �                     &@        �       �                   xp@�k~X��?1             R@        �       �       	          433�?`2U0*��?             9@        �       �                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �        !            �G@        �       �                    �?�q��/��?#            �H@       �       �                    �?r�q��?             B@        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �?��hJ,�?             A@       �       �                   �Z@��a�n`�?             ?@        �       �                   0a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?h�����?             <@        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                   �]@�q�q�?             @        ������������������������       �                     �?        �       �                    �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        �       �       	             @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     �?        �       �                    �?>���Rp�?             =@        �       �                   �[@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `c@�z�G��?             4@        ������������������������       �                      @        �       �                   @`@      �?	             (@        ������������������������       �                     @        �       �                   �g@�q�q�?             "@        ������������������������       �                     �?        �       �                    �H@      �?              @        �       �                   e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  6n����?�� ���?��P�z�?�^�
��?l�l��?�'}�'}�?΀Pr��?����6b�?�;����?br1��?              �?UUUUUU�?UUUUUU�?ӛ���7�?d!Y�B�?�������?�������?              �?�q�q�?�q�q�?      �?        �������?UUUUUU�?      �?                      �?      �?        ������?����>�?a���{�?��{a�?      �?        �؉�؉�?��N��N�?�؉�؉�?ى�؉��?              �?      �?      �?      �?                      �?              �?333333�?�������?;�;��?;�;��?      �?      �?      �?                      �?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?۶m۶m�?%I�$I��?��蕱�?5'��Ps�?tl��?J��8D�?      �?        +�3�=l�?��c.��?UUUUUU�?UUUUUU�?              �?      �?        a��"��?�L[���?              �?�]����?6��9�?�z�G��?{�G�z�?=��<���?�a�a�?      �?        �������?�������?      �?                      �?      �?      �?              �?      �?        zӛ����?d!Y�B�?      �?        ��<��<�?�a�a�?      �?        ��y��y�?�a�a�?      �?        UUUUUU�?UUUUUU�?              �?      �?        6��P^C�?(������?      �?        wwwwww�?�?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?1�0��?�y��y��?�������?ZZZZZZ�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        a���{�?��=���?�������?�������?      �?                      �?              �?      �?      �?      �?              �?      �?      �?                      �?�������?�:��:��?              �?C��6�S�?ާ�d��?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?�m۶m��?�$I�$I�?t�E]t�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?333333�?�������?              �?      �?              �?        ������?�P^Cy�?F]t�E�?]t�E�?      �?      �?�E]t��?]t�E]�?              �?      �?      �?      �?        �������?�������?              �?      �?                      �?;����?|��r��?"pc�
�?��i�V��?�n�Տ?�GJȩ��?              �?�?�������?      �?        ��k���?1P�M��?              �?�q�q�?�8��8��?{�G�z�?���Q��?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?և���X�?/����?UUUUUU�?�������?      �?      �?      �?                      �?�������?KKKKKK�?�c�1Ƹ?�s�9��?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �i��F�?GX�i���?�q�q�?�q�q�?              �?      �?        ffffff�?333333�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�BHzhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKͅ�h��B@3         \       	          ����?�[��N�?�           ��@               !       
             �?��)��?�            �v@                                  �_@��>4��?H             \@                      	          hff�? pƵHP�?#             J@       ������������������������       �                    �G@                                  �\@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        	                           pq@�z�G��?%             N@       
              	          ����?�û��|�?             G@                                  @z�G�z�?             9@                                  �\@      �?             $@        ������������������������       �                      @                                  �h@      �?              @        ������������������������       �                      @                                   �?r�q��?             @       ������������������������       �                     @                                  �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@                                   �?�ՙ/�?             5@        ������������������������       �                     @                                   �?և���X�?	             ,@        ������������������������       �                     @                                  �m@z�G�z�?             $@                                 �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        "       A                    �?0�|#�p�?�            �o@       #       :                    �?�R�+�0�?b            `e@       $       +                   @n@�;u�,a�?Y            �c@       %       &                    @���1��?8            �Z@       ������������������������       �        ,             U@        '       *                     G@�nkK�?             7@        (       )                   @^@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             3@        ,       9                   0d@�:�]��?!            �I@       -       0                   @[@�r����?             >@        .       /                   �c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        1       2                    �?$�q-�?             :@        ������������������������       �                     &@        3       4                   hp@�r����?	             .@        ������������������������       �                     �?        5       6                    �M@@4և���?             ,@       ������������������������       �                     $@        7       8                   �t@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        ;       <                    @�n_Y�K�?	             *@       ������������������������       �                     @        =       >       	          ,33ӿ����X�?             @        ������������������������       �                      @        ?       @                    ]@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        B       Y                    �?��s����?1             U@       C       L                    @�S����?-             S@       D       I                    �?�>����?              K@       E       F                   �p@`Jj��?             ?@       ������������������������       �                     <@        G       H                   (u@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        J       K                    T@���}<S�?             7@        ������������������������       �                      @        ������������������������       �                     5@        M       R                     K@���|���?             6@       N       Q                    �F@8�Z$���?             *@        O       P                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        S       X                   p`@�q�q�?             "@       T       U                   @Y@؇���X�?             @        ������������������������       �                     @        V       W                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        Z       [                     @      �?              @        ������������������������       �                     @        ������������������������       �                     @        ]       �                    �?ByL5���?�            �v@        ^       �                   �r@������?M            �[@       _       �                    �P@r֛w���?B            @W@       `       y                    @R���Q�?:             T@        a       r       	             @X�<ݚ�?             B@       b       e                    �?��
ц��?             :@        c       d                   Xq@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        f       g                    ^@�����?             3@        ������������������������       �                      @        h       k       	          ����?������?             1@        i       j                   `b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       q                   d@؇���X�?             ,@       m       p                   �c@�<ݚ�?             "@       n       o                   Pf@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        s       t                   �]@z�G�z�?             $@        ������������������������       �                     �?        u       v                    �?�����H�?             "@       ������������������������       �                     @        w       x                    \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        z       �       
             �?���7�?             F@       {       |                    �? ���J��?            �C@        ������������������������       �                     6@        }       �                    `@�IєX�?             1@        ~              
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        �       �       	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          033�?��
ц��?             *@        ������������������������       �                     @        �       �                    �?�z�G��?             $@        ������������������������       �                      @        �       �                   @]@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �s@�����H�?             2@        ������������������������       �                     @        �       �       	          ����?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        �       �                    �?     ��?�             p@        �       �                   �f@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?�-���e�?�            �o@       �       �                    @��8"W�?�            �l@        �       �                   �a@R���Q�?             D@       ������������������������       �                     3@        �       �       	          ����?����X�?	             5@        �       �                    �?�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �L@���N8�?z            �g@       �       �                    �?���l��?H            �[@       �       �       
             �?���}<S�?:             W@        ������������������������       �                      @        �       �                   ``@�����?6             U@       �       �                   0f@&^�)b�?            �E@        ������������������������       �                     $@        �       �                   �a@r٣����?            �@@       �       �                   `i@l��
I��?             ;@        �       �                    �E@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �`@��<b���?             7@       �       �                   �s@"pc�
�?             6@       �       �       	          ���@R���Q�?             4@       �       �                     L@�IєX�?
             1@       ������������������������       �        	             0@        ������������������������       �                     �?        �       �                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        ������������������������       �                     3@        �       �       	          ����?�(�Tw�?2            �S@        �       �                     O@�C��2(�?	             &@        �       �                     N@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        )            �P@        �       �                   �_@8����?             7@        ������������������������       �                     "@        �       �                   �`@      �?             ,@       �       �                    �?�<ݚ�?             "@       �       �       	          033�?      �?              @        �       �       	          033�?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  B~�9�J�?�@c�Z�?Np	���?d����?n۶m۶�?%I�$I��?;�;��?'vb'vb�?              �?�������?�������?              �?      �?        333333�?ffffff�?��,d!�?8��Moz�?�������?�������?      �?      �?              �?      �?      �?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?�<��<��?�a�a�?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?      �?      �?      �?                      �?      �?      �?              �?      �?                      �?�������?�?�;�� �?�A|�?�]-n���?h *�3�?�S�rp��?�+J�#�?      �?        �Mozӛ�?d!Y�B�?      �?      �?      �?                      �?      �?        }}}}}}�?�?�������?�?      �?      �?              �?      �?        �؉�؉�?;�;��?      �?        �������?�?              �?n۶m۶�?�$I�$I�?      �?              �?      �?      �?                      �?      �?        ;�;��?ى�؉��?      �?        �$I�$I�?�m۶m��?              �?�������?333333�?              �?      �?        z��y���?�a�a�?(������?^Cy�5�?�Kh/��?h/�����?���{��?�B!��?      �?        UUUUUU�?UUUUUU�?              �?      �?        ӛ���7�?d!Y�B�?              �?      �?        ]t�E]�?F]t�E�?;�;��?;�;��?333333�?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?�7PØ��?�+�U�?q��$�?G���w�?�B!��?���{��?�������?�������?�q�q�?r�q��?�;�;�?�؉�؉�?�$I�$I�?۶m۶m�?              �?      �?        Q^Cy��?^Cy�5�?              �?xxxxxx�?�?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?9��8���?�q�q�?      �?      �?              �?      �?                      �?      �?        �������?�������?      �?        �q�q�?�q�q�?              �?      �?      �?      �?                      �?F]t�E�?�.�袋�?�A�A�?��-��-�?              �?�?�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?                      �?�؉�؉�?�;�;�?      �?        333333�?ffffff�?      �?              �?      �?      �?                      �?�q�q�?�q�q�?      �?        /�袋.�?F]t�E�?      �?                      �?      �?     ��?      �?      �?      �?                      �?�eY�eY�?M�4M�4�?�G�İ?b��g��?333333�?333333�?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?�a�a�?��y��y�?5'��Ps�?��蕱�?d!Y�B�?ӛ���7�?              �?�a�a�?=��<���?�}A_��?���/��?              �?|���?>���>�?h/�����?Lh/����?      �?      �?              �?      �?        ��Moz��?��,d!�?F]t�E�?/�袋.�?333333�?333333�?�?�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?              �?                      �?              �?              �?�A�A�?p��o���?F]t�E�?]t�E�?      �?      �?              �?      �?      �?      �?                      �?              �?              �?8��Moz�?d!Y�B�?              �?      �?      �?9��8���?�q�q�?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?�t�bubhhubehhub.